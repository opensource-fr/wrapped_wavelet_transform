magic
tech sky130A
magscale 1 2
timestamp 1654486978
<< obsli1 >>
rect 1104 2159 58880 57681
<< obsm1 >>
rect 382 1980 59326 58132
<< metal2 >>
rect 634 59200 746 60000
rect 1278 59200 1390 60000
rect 2566 59200 2678 60000
rect 3854 59200 3966 60000
rect 5142 59200 5254 60000
rect 5786 59200 5898 60000
rect 7074 59200 7186 60000
rect 8362 59200 8474 60000
rect 9650 59200 9762 60000
rect 10294 59200 10406 60000
rect 11582 59200 11694 60000
rect 12870 59200 12982 60000
rect 13514 59200 13626 60000
rect 14802 59200 14914 60000
rect 16090 59200 16202 60000
rect 17378 59200 17490 60000
rect 18022 59200 18134 60000
rect 19310 59200 19422 60000
rect 20598 59200 20710 60000
rect 21242 59200 21354 60000
rect 22530 59200 22642 60000
rect 23818 59200 23930 60000
rect 25106 59200 25218 60000
rect 25750 59200 25862 60000
rect 27038 59200 27150 60000
rect 28326 59200 28438 60000
rect 28970 59200 29082 60000
rect 30258 59200 30370 60000
rect 31546 59200 31658 60000
rect 32834 59200 32946 60000
rect 33478 59200 33590 60000
rect 34766 59200 34878 60000
rect 36054 59200 36166 60000
rect 36698 59200 36810 60000
rect 37986 59200 38098 60000
rect 39274 59200 39386 60000
rect 40562 59200 40674 60000
rect 41206 59200 41318 60000
rect 42494 59200 42606 60000
rect 43782 59200 43894 60000
rect 44426 59200 44538 60000
rect 45714 59200 45826 60000
rect 47002 59200 47114 60000
rect 48290 59200 48402 60000
rect 48934 59200 49046 60000
rect 50222 59200 50334 60000
rect 51510 59200 51622 60000
rect 52154 59200 52266 60000
rect 53442 59200 53554 60000
rect 54730 59200 54842 60000
rect 56018 59200 56130 60000
rect 56662 59200 56774 60000
rect 57950 59200 58062 60000
rect 59238 59200 59350 60000
rect 59882 59200 59994 60000
rect -10 0 102 800
rect 634 0 746 800
rect 1922 0 2034 800
rect 3210 0 3322 800
rect 3854 0 3966 800
rect 5142 0 5254 800
rect 6430 0 6542 800
rect 7718 0 7830 800
rect 8362 0 8474 800
rect 9650 0 9762 800
rect 10938 0 11050 800
rect 11582 0 11694 800
rect 12870 0 12982 800
rect 14158 0 14270 800
rect 15446 0 15558 800
rect 16090 0 16202 800
rect 17378 0 17490 800
rect 18666 0 18778 800
rect 19310 0 19422 800
rect 20598 0 20710 800
rect 21886 0 21998 800
rect 23174 0 23286 800
rect 23818 0 23930 800
rect 25106 0 25218 800
rect 26394 0 26506 800
rect 27038 0 27150 800
rect 28326 0 28438 800
rect 29614 0 29726 800
rect 30902 0 31014 800
rect 31546 0 31658 800
rect 32834 0 32946 800
rect 34122 0 34234 800
rect 34766 0 34878 800
rect 36054 0 36166 800
rect 37342 0 37454 800
rect 38630 0 38742 800
rect 39274 0 39386 800
rect 40562 0 40674 800
rect 41850 0 41962 800
rect 42494 0 42606 800
rect 43782 0 43894 800
rect 45070 0 45182 800
rect 46358 0 46470 800
rect 47002 0 47114 800
rect 48290 0 48402 800
rect 49578 0 49690 800
rect 50222 0 50334 800
rect 51510 0 51622 800
rect 52798 0 52910 800
rect 54086 0 54198 800
rect 54730 0 54842 800
rect 56018 0 56130 800
rect 57306 0 57418 800
rect 58594 0 58706 800
rect 59238 0 59350 800
<< obsm2 >>
rect 386 59144 578 59200
rect 802 59144 1222 59200
rect 1446 59144 2510 59200
rect 2734 59144 3798 59200
rect 4022 59144 5086 59200
rect 5310 59144 5730 59200
rect 5954 59144 7018 59200
rect 7242 59144 8306 59200
rect 8530 59144 9594 59200
rect 9818 59144 10238 59200
rect 10462 59144 11526 59200
rect 11750 59144 12814 59200
rect 13038 59144 13458 59200
rect 13682 59144 14746 59200
rect 14970 59144 16034 59200
rect 16258 59144 17322 59200
rect 17546 59144 17966 59200
rect 18190 59144 19254 59200
rect 19478 59144 20542 59200
rect 20766 59144 21186 59200
rect 21410 59144 22474 59200
rect 22698 59144 23762 59200
rect 23986 59144 25050 59200
rect 25274 59144 25694 59200
rect 25918 59144 26982 59200
rect 27206 59144 28270 59200
rect 28494 59144 28914 59200
rect 29138 59144 30202 59200
rect 30426 59144 31490 59200
rect 31714 59144 32778 59200
rect 33002 59144 33422 59200
rect 33646 59144 34710 59200
rect 34934 59144 35998 59200
rect 36222 59144 36642 59200
rect 36866 59144 37930 59200
rect 38154 59144 39218 59200
rect 39442 59144 40506 59200
rect 40730 59144 41150 59200
rect 41374 59144 42438 59200
rect 42662 59144 43726 59200
rect 43950 59144 44370 59200
rect 44594 59144 45658 59200
rect 45882 59144 46946 59200
rect 47170 59144 48234 59200
rect 48458 59144 48878 59200
rect 49102 59144 50166 59200
rect 50390 59144 51454 59200
rect 51678 59144 52098 59200
rect 52322 59144 53386 59200
rect 53610 59144 54674 59200
rect 54898 59144 55962 59200
rect 56186 59144 56606 59200
rect 56830 59144 57894 59200
rect 58118 59144 59182 59200
rect 386 856 59320 59144
rect 386 31 578 856
rect 802 31 1866 856
rect 2090 31 3154 856
rect 3378 31 3798 856
rect 4022 31 5086 856
rect 5310 31 6374 856
rect 6598 31 7662 856
rect 7886 31 8306 856
rect 8530 31 9594 856
rect 9818 31 10882 856
rect 11106 31 11526 856
rect 11750 31 12814 856
rect 13038 31 14102 856
rect 14326 31 15390 856
rect 15614 31 16034 856
rect 16258 31 17322 856
rect 17546 31 18610 856
rect 18834 31 19254 856
rect 19478 31 20542 856
rect 20766 31 21830 856
rect 22054 31 23118 856
rect 23342 31 23762 856
rect 23986 31 25050 856
rect 25274 31 26338 856
rect 26562 31 26982 856
rect 27206 31 28270 856
rect 28494 31 29558 856
rect 29782 31 30846 856
rect 31070 31 31490 856
rect 31714 31 32778 856
rect 33002 31 34066 856
rect 34290 31 34710 856
rect 34934 31 35998 856
rect 36222 31 37286 856
rect 37510 31 38574 856
rect 38798 31 39218 856
rect 39442 31 40506 856
rect 40730 31 41794 856
rect 42018 31 42438 856
rect 42662 31 43726 856
rect 43950 31 45014 856
rect 45238 31 46302 856
rect 46526 31 46946 856
rect 47170 31 48234 856
rect 48458 31 49522 856
rect 49746 31 50166 856
rect 50390 31 51454 856
rect 51678 31 52742 856
rect 52966 31 54030 856
rect 54254 31 54674 856
rect 54898 31 55962 856
rect 56186 31 57250 856
rect 57474 31 58538 856
rect 58762 31 59182 856
<< metal3 >>
rect 0 59108 800 59348
rect 59200 58428 60000 58668
rect 0 57748 800 57988
rect 0 57068 800 57308
rect 59200 57068 60000 57308
rect 0 55708 800 55948
rect 59200 55708 60000 55948
rect 59200 55028 60000 55268
rect 0 54348 800 54588
rect 59200 53668 60000 53908
rect 0 52988 800 53228
rect 0 52308 800 52548
rect 59200 52308 60000 52548
rect 0 50948 800 51188
rect 59200 50948 60000 51188
rect 59200 50268 60000 50508
rect 0 49588 800 49828
rect 0 48908 800 49148
rect 59200 48908 60000 49148
rect 0 47548 800 47788
rect 59200 47548 60000 47788
rect 59200 46868 60000 47108
rect 0 46188 800 46428
rect 59200 45508 60000 45748
rect 0 44828 800 45068
rect 0 44148 800 44388
rect 59200 44148 60000 44388
rect 0 42788 800 43028
rect 59200 42788 60000 43028
rect 59200 42108 60000 42348
rect 0 41428 800 41668
rect 0 40748 800 40988
rect 59200 40748 60000 40988
rect 0 39388 800 39628
rect 59200 39388 60000 39628
rect 59200 38708 60000 38948
rect 0 38028 800 38268
rect 59200 37348 60000 37588
rect 0 36668 800 36908
rect 0 35988 800 36228
rect 59200 35988 60000 36228
rect 0 34628 800 34868
rect 59200 34628 60000 34868
rect 59200 33948 60000 34188
rect 0 33268 800 33508
rect 0 32588 800 32828
rect 59200 32588 60000 32828
rect 0 31228 800 31468
rect 59200 31228 60000 31468
rect 59200 30548 60000 30788
rect 0 29868 800 30108
rect 59200 29188 60000 29428
rect 0 28508 800 28748
rect 0 27828 800 28068
rect 59200 27828 60000 28068
rect 0 26468 800 26708
rect 59200 26468 60000 26708
rect 59200 25788 60000 26028
rect 0 25108 800 25348
rect 0 24428 800 24668
rect 59200 24428 60000 24668
rect 0 23068 800 23308
rect 59200 23068 60000 23308
rect 59200 22388 60000 22628
rect 0 21708 800 21948
rect 59200 21028 60000 21268
rect 0 20348 800 20588
rect 0 19668 800 19908
rect 59200 19668 60000 19908
rect 0 18308 800 18548
rect 59200 18308 60000 18548
rect 59200 17628 60000 17868
rect 0 16948 800 17188
rect 0 16268 800 16508
rect 59200 16268 60000 16508
rect 0 14908 800 15148
rect 59200 14908 60000 15148
rect 59200 14228 60000 14468
rect 0 13548 800 13788
rect 59200 12868 60000 13108
rect 0 12188 800 12428
rect 0 11508 800 11748
rect 59200 11508 60000 11748
rect 0 10148 800 10388
rect 59200 10148 60000 10388
rect 59200 9468 60000 9708
rect 0 8788 800 9028
rect 0 8108 800 8348
rect 59200 8108 60000 8348
rect 0 6748 800 6988
rect 59200 6748 60000 6988
rect 59200 6068 60000 6308
rect 0 5388 800 5628
rect 59200 4708 60000 4948
rect 0 4028 800 4268
rect 0 3348 800 3588
rect 59200 3348 60000 3588
rect 0 1988 800 2228
rect 59200 1988 60000 2228
rect 59200 1308 60000 1548
rect 0 628 800 868
rect 59200 -52 60000 188
<< obsm3 >>
rect 381 58348 59120 58581
rect 381 58068 59235 58348
rect 880 57668 59235 58068
rect 381 57388 59235 57668
rect 880 56988 59120 57388
rect 381 56028 59235 56988
rect 880 55628 59120 56028
rect 381 55348 59235 55628
rect 381 54948 59120 55348
rect 381 54668 59235 54948
rect 880 54268 59235 54668
rect 381 53988 59235 54268
rect 381 53588 59120 53988
rect 381 53308 59235 53588
rect 880 52908 59235 53308
rect 381 52628 59235 52908
rect 880 52228 59120 52628
rect 381 51268 59235 52228
rect 880 50868 59120 51268
rect 381 50588 59235 50868
rect 381 50188 59120 50588
rect 381 49908 59235 50188
rect 880 49508 59235 49908
rect 381 49228 59235 49508
rect 880 48828 59120 49228
rect 381 47868 59235 48828
rect 880 47468 59120 47868
rect 381 47188 59235 47468
rect 381 46788 59120 47188
rect 381 46508 59235 46788
rect 880 46108 59235 46508
rect 381 45828 59235 46108
rect 381 45428 59120 45828
rect 381 45148 59235 45428
rect 880 44748 59235 45148
rect 381 44468 59235 44748
rect 880 44068 59120 44468
rect 381 43108 59235 44068
rect 880 42708 59120 43108
rect 381 42428 59235 42708
rect 381 42028 59120 42428
rect 381 41748 59235 42028
rect 880 41348 59235 41748
rect 381 41068 59235 41348
rect 880 40668 59120 41068
rect 381 39708 59235 40668
rect 880 39308 59120 39708
rect 381 39028 59235 39308
rect 381 38628 59120 39028
rect 381 38348 59235 38628
rect 880 37948 59235 38348
rect 381 37668 59235 37948
rect 381 37268 59120 37668
rect 381 36988 59235 37268
rect 880 36588 59235 36988
rect 381 36308 59235 36588
rect 880 35908 59120 36308
rect 381 34948 59235 35908
rect 880 34548 59120 34948
rect 381 34268 59235 34548
rect 381 33868 59120 34268
rect 381 33588 59235 33868
rect 880 33188 59235 33588
rect 381 32908 59235 33188
rect 880 32508 59120 32908
rect 381 31548 59235 32508
rect 880 31148 59120 31548
rect 381 30868 59235 31148
rect 381 30468 59120 30868
rect 381 30188 59235 30468
rect 880 29788 59235 30188
rect 381 29508 59235 29788
rect 381 29108 59120 29508
rect 381 28828 59235 29108
rect 880 28428 59235 28828
rect 381 28148 59235 28428
rect 880 27748 59120 28148
rect 381 26788 59235 27748
rect 880 26388 59120 26788
rect 381 26108 59235 26388
rect 381 25708 59120 26108
rect 381 25428 59235 25708
rect 880 25028 59235 25428
rect 381 24748 59235 25028
rect 880 24348 59120 24748
rect 381 23388 59235 24348
rect 880 22988 59120 23388
rect 381 22708 59235 22988
rect 381 22308 59120 22708
rect 381 22028 59235 22308
rect 880 21628 59235 22028
rect 381 21348 59235 21628
rect 381 20948 59120 21348
rect 381 20668 59235 20948
rect 880 20268 59235 20668
rect 381 19988 59235 20268
rect 880 19588 59120 19988
rect 381 18628 59235 19588
rect 880 18228 59120 18628
rect 381 17948 59235 18228
rect 381 17548 59120 17948
rect 381 17268 59235 17548
rect 880 16868 59235 17268
rect 381 16588 59235 16868
rect 880 16188 59120 16588
rect 381 15228 59235 16188
rect 880 14828 59120 15228
rect 381 14548 59235 14828
rect 381 14148 59120 14548
rect 381 13868 59235 14148
rect 880 13468 59235 13868
rect 381 13188 59235 13468
rect 381 12788 59120 13188
rect 381 12508 59235 12788
rect 880 12108 59235 12508
rect 381 11828 59235 12108
rect 880 11428 59120 11828
rect 381 10468 59235 11428
rect 880 10068 59120 10468
rect 381 9788 59235 10068
rect 381 9388 59120 9788
rect 381 9108 59235 9388
rect 880 8708 59235 9108
rect 381 8428 59235 8708
rect 880 8028 59120 8428
rect 381 7068 59235 8028
rect 880 6668 59120 7068
rect 381 6388 59235 6668
rect 381 5988 59120 6388
rect 381 5708 59235 5988
rect 880 5308 59235 5708
rect 381 5028 59235 5308
rect 381 4628 59120 5028
rect 381 4348 59235 4628
rect 880 3948 59235 4348
rect 381 3668 59235 3948
rect 880 3268 59120 3668
rect 381 2308 59235 3268
rect 880 1908 59120 2308
rect 381 1628 59235 1908
rect 381 1228 59120 1628
rect 381 948 59235 1228
rect 880 548 59235 948
rect 381 268 59235 548
rect 381 35 59120 268
<< metal4 >>
rect 4208 2128 4528 57712
rect 19568 2128 19888 57712
rect 34928 2128 35248 57712
rect 50288 2128 50608 57712
<< obsm4 >>
rect 1899 5747 4128 57629
rect 4608 5747 19488 57629
rect 19968 5747 34848 57629
rect 35328 5747 50208 57629
rect 50688 5747 57717 57629
<< labels >>
rlabel metal3 s 0 55708 800 55948 6 active
port 1 nsew signal input
rlabel metal2 s 18666 0 18778 800 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 33478 59200 33590 60000 6 io_in[10]
port 3 nsew signal input
rlabel metal2 s 634 59200 746 60000 6 io_in[11]
port 4 nsew signal input
rlabel metal3 s 59200 50268 60000 50508 6 io_in[12]
port 5 nsew signal input
rlabel metal2 s 28326 0 28438 800 6 io_in[13]
port 6 nsew signal input
rlabel metal2 s 22530 59200 22642 60000 6 io_in[14]
port 7 nsew signal input
rlabel metal3 s 59200 52308 60000 52548 6 io_in[15]
port 8 nsew signal input
rlabel metal3 s 59200 4708 60000 4948 6 io_in[16]
port 9 nsew signal input
rlabel metal2 s 12870 59200 12982 60000 6 io_in[17]
port 10 nsew signal input
rlabel metal2 s 14802 59200 14914 60000 6 io_in[18]
port 11 nsew signal input
rlabel metal2 s 51510 0 51622 800 6 io_in[19]
port 12 nsew signal input
rlabel metal3 s 0 19668 800 19908 6 io_in[1]
port 13 nsew signal input
rlabel metal3 s 0 34628 800 34868 6 io_in[20]
port 14 nsew signal input
rlabel metal3 s 0 23068 800 23308 6 io_in[21]
port 15 nsew signal input
rlabel metal3 s 59200 18308 60000 18548 6 io_in[22]
port 16 nsew signal input
rlabel metal2 s 11582 59200 11694 60000 6 io_in[23]
port 17 nsew signal input
rlabel metal2 s 8362 59200 8474 60000 6 io_in[24]
port 18 nsew signal input
rlabel metal2 s 45070 0 45182 800 6 io_in[25]
port 19 nsew signal input
rlabel metal2 s 43782 0 43894 800 6 io_in[26]
port 20 nsew signal input
rlabel metal3 s 59200 12868 60000 13108 6 io_in[27]
port 21 nsew signal input
rlabel metal2 s 39274 0 39386 800 6 io_in[28]
port 22 nsew signal input
rlabel metal2 s 59882 59200 59994 60000 6 io_in[29]
port 23 nsew signal input
rlabel metal2 s 19310 0 19422 800 6 io_in[2]
port 24 nsew signal input
rlabel metal3 s 59200 23068 60000 23308 6 io_in[30]
port 25 nsew signal input
rlabel metal3 s 0 52988 800 53228 6 io_in[31]
port 26 nsew signal input
rlabel metal2 s 37342 0 37454 800 6 io_in[32]
port 27 nsew signal input
rlabel metal3 s 0 31228 800 31468 6 io_in[33]
port 28 nsew signal input
rlabel metal2 s 45714 59200 45826 60000 6 io_in[34]
port 29 nsew signal input
rlabel metal2 s 52154 59200 52266 60000 6 io_in[35]
port 30 nsew signal input
rlabel metal3 s 59200 37348 60000 37588 6 io_in[36]
port 31 nsew signal input
rlabel metal2 s 53442 59200 53554 60000 6 io_in[37]
port 32 nsew signal input
rlabel metal2 s 34766 59200 34878 60000 6 io_in[3]
port 33 nsew signal input
rlabel metal3 s 59200 35988 60000 36228 6 io_in[4]
port 34 nsew signal input
rlabel metal3 s 59200 57068 60000 57308 6 io_in[5]
port 35 nsew signal input
rlabel metal3 s 0 36668 800 36908 6 io_in[6]
port 36 nsew signal input
rlabel metal3 s 0 25108 800 25348 6 io_in[7]
port 37 nsew signal input
rlabel metal3 s 59200 39388 60000 39628 6 io_in[8]
port 38 nsew signal input
rlabel metal2 s 10294 59200 10406 60000 6 io_in[9]
port 39 nsew signal input
rlabel metal2 s 31546 0 31658 800 6 io_oeb[0]
port 40 nsew signal bidirectional
rlabel metal3 s 0 20348 800 20588 6 io_oeb[10]
port 41 nsew signal bidirectional
rlabel metal3 s 59200 33948 60000 34188 6 io_oeb[11]
port 42 nsew signal bidirectional
rlabel metal3 s 59200 17628 60000 17868 6 io_oeb[12]
port 43 nsew signal bidirectional
rlabel metal3 s 59200 16268 60000 16508 6 io_oeb[13]
port 44 nsew signal bidirectional
rlabel metal3 s 0 5388 800 5628 6 io_oeb[14]
port 45 nsew signal bidirectional
rlabel metal2 s 17378 59200 17490 60000 6 io_oeb[15]
port 46 nsew signal bidirectional
rlabel metal3 s 59200 1988 60000 2228 6 io_oeb[16]
port 47 nsew signal bidirectional
rlabel metal2 s 16090 0 16202 800 6 io_oeb[17]
port 48 nsew signal bidirectional
rlabel metal2 s 43782 59200 43894 60000 6 io_oeb[18]
port 49 nsew signal bidirectional
rlabel metal2 s 18022 59200 18134 60000 6 io_oeb[19]
port 50 nsew signal bidirectional
rlabel metal2 s 47002 0 47114 800 6 io_oeb[1]
port 51 nsew signal bidirectional
rlabel metal3 s 59200 25788 60000 26028 6 io_oeb[20]
port 52 nsew signal bidirectional
rlabel metal2 s 2566 59200 2678 60000 6 io_oeb[21]
port 53 nsew signal bidirectional
rlabel metal2 s 6430 0 6542 800 6 io_oeb[22]
port 54 nsew signal bidirectional
rlabel metal2 s 30258 59200 30370 60000 6 io_oeb[23]
port 55 nsew signal bidirectional
rlabel metal2 s 31546 59200 31658 60000 6 io_oeb[24]
port 56 nsew signal bidirectional
rlabel metal2 s 57306 0 57418 800 6 io_oeb[25]
port 57 nsew signal bidirectional
rlabel metal3 s 59200 46868 60000 47108 6 io_oeb[26]
port 58 nsew signal bidirectional
rlabel metal2 s 36054 59200 36166 60000 6 io_oeb[27]
port 59 nsew signal bidirectional
rlabel metal2 s 50222 0 50334 800 6 io_oeb[28]
port 60 nsew signal bidirectional
rlabel metal3 s 59200 38708 60000 38948 6 io_oeb[29]
port 61 nsew signal bidirectional
rlabel metal2 s 50222 59200 50334 60000 6 io_oeb[2]
port 62 nsew signal bidirectional
rlabel metal2 s 3854 59200 3966 60000 6 io_oeb[30]
port 63 nsew signal bidirectional
rlabel metal2 s 49578 0 49690 800 6 io_oeb[31]
port 64 nsew signal bidirectional
rlabel metal3 s 0 29868 800 30108 6 io_oeb[32]
port 65 nsew signal bidirectional
rlabel metal2 s 58594 0 58706 800 6 io_oeb[33]
port 66 nsew signal bidirectional
rlabel metal2 s 13514 59200 13626 60000 6 io_oeb[34]
port 67 nsew signal bidirectional
rlabel metal3 s 0 26468 800 26708 6 io_oeb[35]
port 68 nsew signal bidirectional
rlabel metal3 s 0 13548 800 13788 6 io_oeb[36]
port 69 nsew signal bidirectional
rlabel metal3 s 0 21708 800 21948 6 io_oeb[37]
port 70 nsew signal bidirectional
rlabel metal2 s 30902 0 31014 800 6 io_oeb[3]
port 71 nsew signal bidirectional
rlabel metal3 s 59200 -52 60000 188 6 io_oeb[4]
port 72 nsew signal bidirectional
rlabel metal3 s 0 39388 800 39628 6 io_oeb[5]
port 73 nsew signal bidirectional
rlabel metal3 s 59200 21028 60000 21268 6 io_oeb[6]
port 74 nsew signal bidirectional
rlabel metal2 s 16090 59200 16202 60000 6 io_oeb[7]
port 75 nsew signal bidirectional
rlabel metal2 s 5142 0 5254 800 6 io_oeb[8]
port 76 nsew signal bidirectional
rlabel metal2 s 12870 0 12982 800 6 io_oeb[9]
port 77 nsew signal bidirectional
rlabel metal3 s 59200 55708 60000 55948 6 io_out[0]
port 78 nsew signal bidirectional
rlabel metal3 s 59200 32588 60000 32828 6 io_out[10]
port 79 nsew signal bidirectional
rlabel metal3 s 0 3348 800 3588 6 io_out[11]
port 80 nsew signal bidirectional
rlabel metal3 s 0 8788 800 9028 6 io_out[12]
port 81 nsew signal bidirectional
rlabel metal2 s 48290 0 48402 800 6 io_out[13]
port 82 nsew signal bidirectional
rlabel metal3 s 59200 47548 60000 47788 6 io_out[14]
port 83 nsew signal bidirectional
rlabel metal3 s 0 49588 800 49828 6 io_out[15]
port 84 nsew signal bidirectional
rlabel metal3 s 59200 31228 60000 31468 6 io_out[16]
port 85 nsew signal bidirectional
rlabel metal2 s 56018 59200 56130 60000 6 io_out[17]
port 86 nsew signal bidirectional
rlabel metal2 s 56018 0 56130 800 6 io_out[18]
port 87 nsew signal bidirectional
rlabel metal3 s 0 28508 800 28748 6 io_out[19]
port 88 nsew signal bidirectional
rlabel metal2 s 40562 59200 40674 60000 6 io_out[1]
port 89 nsew signal bidirectional
rlabel metal2 s 48934 59200 49046 60000 6 io_out[20]
port 90 nsew signal bidirectional
rlabel metal3 s 0 48908 800 49148 6 io_out[21]
port 91 nsew signal bidirectional
rlabel metal2 s 38630 0 38742 800 6 io_out[22]
port 92 nsew signal bidirectional
rlabel metal3 s 59200 26468 60000 26708 6 io_out[23]
port 93 nsew signal bidirectional
rlabel metal2 s 32834 0 32946 800 6 io_out[24]
port 94 nsew signal bidirectional
rlabel metal2 s 44426 59200 44538 60000 6 io_out[25]
port 95 nsew signal bidirectional
rlabel metal3 s 0 6748 800 6988 6 io_out[26]
port 96 nsew signal bidirectional
rlabel metal2 s 47002 59200 47114 60000 6 io_out[27]
port 97 nsew signal bidirectional
rlabel metal2 s 20598 0 20710 800 6 io_out[28]
port 98 nsew signal bidirectional
rlabel metal3 s 59200 1308 60000 1548 6 io_out[29]
port 99 nsew signal bidirectional
rlabel metal2 s 8362 0 8474 800 6 io_out[2]
port 100 nsew signal bidirectional
rlabel metal3 s 0 8108 800 8348 6 io_out[30]
port 101 nsew signal bidirectional
rlabel metal3 s 0 16948 800 17188 6 io_out[31]
port 102 nsew signal bidirectional
rlabel metal3 s 0 57068 800 57308 6 io_out[32]
port 103 nsew signal bidirectional
rlabel metal3 s 59200 8108 60000 8348 6 io_out[33]
port 104 nsew signal bidirectional
rlabel metal3 s 59200 48908 60000 49148 6 io_out[34]
port 105 nsew signal bidirectional
rlabel metal3 s 59200 45508 60000 45748 6 io_out[35]
port 106 nsew signal bidirectional
rlabel metal2 s 19310 59200 19422 60000 6 io_out[36]
port 107 nsew signal bidirectional
rlabel metal3 s 59200 53668 60000 53908 6 io_out[37]
port 108 nsew signal bidirectional
rlabel metal3 s 0 52308 800 52548 6 io_out[3]
port 109 nsew signal bidirectional
rlabel metal3 s 59200 34628 60000 34868 6 io_out[4]
port 110 nsew signal bidirectional
rlabel metal2 s 28326 59200 28438 60000 6 io_out[5]
port 111 nsew signal bidirectional
rlabel metal2 s 57950 59200 58062 60000 6 io_out[6]
port 112 nsew signal bidirectional
rlabel metal3 s 0 24428 800 24668 6 io_out[7]
port 113 nsew signal bidirectional
rlabel metal2 s 23174 0 23286 800 6 io_out[8]
port 114 nsew signal bidirectional
rlabel metal3 s 0 18308 800 18548 6 io_out[9]
port 115 nsew signal bidirectional
rlabel metal3 s 59200 9468 60000 9708 6 la1_data_in[0]
port 116 nsew signal input
rlabel metal2 s 26394 0 26506 800 6 la1_data_in[10]
port 117 nsew signal input
rlabel metal3 s 59200 6748 60000 6988 6 la1_data_in[11]
port 118 nsew signal input
rlabel metal3 s 0 44828 800 45068 6 la1_data_in[12]
port 119 nsew signal input
rlabel metal2 s 40562 0 40674 800 6 la1_data_in[13]
port 120 nsew signal input
rlabel metal3 s 0 16268 800 16508 6 la1_data_in[14]
port 121 nsew signal input
rlabel metal2 s 20598 59200 20710 60000 6 la1_data_in[15]
port 122 nsew signal input
rlabel metal2 s 37986 59200 38098 60000 6 la1_data_in[16]
port 123 nsew signal input
rlabel metal2 s 28970 59200 29082 60000 6 la1_data_in[17]
port 124 nsew signal input
rlabel metal2 s 52798 0 52910 800 6 la1_data_in[18]
port 125 nsew signal input
rlabel metal2 s 21242 59200 21354 60000 6 la1_data_in[19]
port 126 nsew signal input
rlabel metal2 s 23818 0 23930 800 6 la1_data_in[1]
port 127 nsew signal input
rlabel metal3 s 0 44148 800 44388 6 la1_data_in[20]
port 128 nsew signal input
rlabel metal2 s 59238 59200 59350 60000 6 la1_data_in[21]
port 129 nsew signal input
rlabel metal3 s 59200 10148 60000 10388 6 la1_data_in[22]
port 130 nsew signal input
rlabel metal3 s 0 628 800 868 6 la1_data_in[23]
port 131 nsew signal input
rlabel metal2 s 17378 0 17490 800 6 la1_data_in[24]
port 132 nsew signal input
rlabel metal3 s 0 46188 800 46428 6 la1_data_in[25]
port 133 nsew signal input
rlabel metal3 s 59200 3348 60000 3588 6 la1_data_in[26]
port 134 nsew signal input
rlabel metal2 s 34766 0 34878 800 6 la1_data_in[27]
port 135 nsew signal input
rlabel metal3 s 0 40748 800 40988 6 la1_data_in[28]
port 136 nsew signal input
rlabel metal2 s 1278 59200 1390 60000 6 la1_data_in[29]
port 137 nsew signal input
rlabel metal2 s 14158 0 14270 800 6 la1_data_in[2]
port 138 nsew signal input
rlabel metal2 s 1922 0 2034 800 6 la1_data_in[30]
port 139 nsew signal input
rlabel metal2 s 46358 0 46470 800 6 la1_data_in[31]
port 140 nsew signal input
rlabel metal3 s 0 38028 800 38268 6 la1_data_in[3]
port 141 nsew signal input
rlabel metal2 s 51510 59200 51622 60000 6 la1_data_in[4]
port 142 nsew signal input
rlabel metal3 s 59200 29188 60000 29428 6 la1_data_in[5]
port 143 nsew signal input
rlabel metal2 s 23818 59200 23930 60000 6 la1_data_in[6]
port 144 nsew signal input
rlabel metal3 s 0 27828 800 28068 6 la1_data_in[7]
port 145 nsew signal input
rlabel metal2 s 25106 59200 25218 60000 6 la1_data_in[8]
port 146 nsew signal input
rlabel metal3 s 0 41428 800 41668 6 la1_data_in[9]
port 147 nsew signal input
rlabel metal2 s 9650 0 9762 800 6 la1_data_out[0]
port 148 nsew signal bidirectional
rlabel metal3 s 59200 14228 60000 14468 6 la1_data_out[10]
port 149 nsew signal bidirectional
rlabel metal2 s 27038 0 27150 800 6 la1_data_out[11]
port 150 nsew signal bidirectional
rlabel metal3 s 59200 55028 60000 55268 6 la1_data_out[12]
port 151 nsew signal bidirectional
rlabel metal2 s 5786 59200 5898 60000 6 la1_data_out[13]
port 152 nsew signal bidirectional
rlabel metal2 s 32834 59200 32946 60000 6 la1_data_out[14]
port 153 nsew signal bidirectional
rlabel metal3 s 0 1988 800 2228 6 la1_data_out[15]
port 154 nsew signal bidirectional
rlabel metal3 s 59200 19668 60000 19908 6 la1_data_out[16]
port 155 nsew signal bidirectional
rlabel metal3 s 59200 42788 60000 43028 6 la1_data_out[17]
port 156 nsew signal bidirectional
rlabel metal2 s 7074 59200 7186 60000 6 la1_data_out[18]
port 157 nsew signal bidirectional
rlabel metal3 s 59200 30548 60000 30788 6 la1_data_out[19]
port 158 nsew signal bidirectional
rlabel metal3 s 0 54348 800 54588 6 la1_data_out[1]
port 159 nsew signal bidirectional
rlabel metal3 s 0 12188 800 12428 6 la1_data_out[20]
port 160 nsew signal bidirectional
rlabel metal3 s 59200 50948 60000 51188 6 la1_data_out[21]
port 161 nsew signal bidirectional
rlabel metal2 s 36698 59200 36810 60000 6 la1_data_out[22]
port 162 nsew signal bidirectional
rlabel metal2 s 15446 0 15558 800 6 la1_data_out[23]
port 163 nsew signal bidirectional
rlabel metal3 s 59200 22388 60000 22628 6 la1_data_out[24]
port 164 nsew signal bidirectional
rlabel metal3 s 0 4028 800 4268 6 la1_data_out[25]
port 165 nsew signal bidirectional
rlabel metal3 s 59200 6068 60000 6308 6 la1_data_out[26]
port 166 nsew signal bidirectional
rlabel metal3 s 0 57748 800 57988 6 la1_data_out[27]
port 167 nsew signal bidirectional
rlabel metal2 s 54086 0 54198 800 6 la1_data_out[28]
port 168 nsew signal bidirectional
rlabel metal2 s 7718 0 7830 800 6 la1_data_out[29]
port 169 nsew signal bidirectional
rlabel metal2 s 25106 0 25218 800 6 la1_data_out[2]
port 170 nsew signal bidirectional
rlabel metal3 s 59200 14908 60000 15148 6 la1_data_out[30]
port 171 nsew signal bidirectional
rlabel metal3 s 59200 58428 60000 58668 6 la1_data_out[31]
port 172 nsew signal bidirectional
rlabel metal3 s 0 11508 800 11748 6 la1_data_out[3]
port 173 nsew signal bidirectional
rlabel metal2 s 54730 0 54842 800 6 la1_data_out[4]
port 174 nsew signal bidirectional
rlabel metal2 s 3854 0 3966 800 6 la1_data_out[5]
port 175 nsew signal bidirectional
rlabel metal3 s 59200 24428 60000 24668 6 la1_data_out[6]
port 176 nsew signal bidirectional
rlabel metal2 s 634 0 746 800 6 la1_data_out[7]
port 177 nsew signal bidirectional
rlabel metal3 s 59200 44148 60000 44388 6 la1_data_out[8]
port 178 nsew signal bidirectional
rlabel metal2 s 56662 59200 56774 60000 6 la1_data_out[9]
port 179 nsew signal bidirectional
rlabel metal2 s 59238 0 59350 800 6 la1_oenb[0]
port 180 nsew signal input
rlabel metal2 s 54730 59200 54842 60000 6 la1_oenb[10]
port 181 nsew signal input
rlabel metal3 s 0 33268 800 33508 6 la1_oenb[11]
port 182 nsew signal input
rlabel metal3 s 0 35988 800 36228 6 la1_oenb[12]
port 183 nsew signal input
rlabel metal2 s 36054 0 36166 800 6 la1_oenb[13]
port 184 nsew signal input
rlabel metal2 s -10 0 102 800 6 la1_oenb[14]
port 185 nsew signal input
rlabel metal2 s 42494 0 42606 800 6 la1_oenb[15]
port 186 nsew signal input
rlabel metal3 s 0 42788 800 43028 6 la1_oenb[16]
port 187 nsew signal input
rlabel metal2 s 5142 59200 5254 60000 6 la1_oenb[17]
port 188 nsew signal input
rlabel metal2 s 27038 59200 27150 60000 6 la1_oenb[18]
port 189 nsew signal input
rlabel metal3 s 0 32588 800 32828 6 la1_oenb[19]
port 190 nsew signal input
rlabel metal2 s 10938 0 11050 800 6 la1_oenb[1]
port 191 nsew signal input
rlabel metal2 s 3210 0 3322 800 6 la1_oenb[20]
port 192 nsew signal input
rlabel metal2 s 39274 59200 39386 60000 6 la1_oenb[21]
port 193 nsew signal input
rlabel metal2 s 25750 59200 25862 60000 6 la1_oenb[22]
port 194 nsew signal input
rlabel metal2 s 29614 0 29726 800 6 la1_oenb[23]
port 195 nsew signal input
rlabel metal2 s 48290 59200 48402 60000 6 la1_oenb[24]
port 196 nsew signal input
rlabel metal3 s 59200 11508 60000 11748 6 la1_oenb[25]
port 197 nsew signal input
rlabel metal3 s 0 47548 800 47788 6 la1_oenb[26]
port 198 nsew signal input
rlabel metal3 s 59200 42108 60000 42348 6 la1_oenb[27]
port 199 nsew signal input
rlabel metal2 s 11582 0 11694 800 6 la1_oenb[28]
port 200 nsew signal input
rlabel metal2 s 21886 0 21998 800 6 la1_oenb[29]
port 201 nsew signal input
rlabel metal3 s 0 10148 800 10388 6 la1_oenb[2]
port 202 nsew signal input
rlabel metal3 s 59200 40748 60000 40988 6 la1_oenb[30]
port 203 nsew signal input
rlabel metal2 s 34122 0 34234 800 6 la1_oenb[31]
port 204 nsew signal input
rlabel metal2 s 42494 59200 42606 60000 6 la1_oenb[3]
port 205 nsew signal input
rlabel metal2 s 41206 59200 41318 60000 6 la1_oenb[4]
port 206 nsew signal input
rlabel metal3 s 0 59108 800 59348 6 la1_oenb[5]
port 207 nsew signal input
rlabel metal2 s 9650 59200 9762 60000 6 la1_oenb[6]
port 208 nsew signal input
rlabel metal2 s 41850 0 41962 800 6 la1_oenb[7]
port 209 nsew signal input
rlabel metal3 s 0 14908 800 15148 6 la1_oenb[8]
port 210 nsew signal input
rlabel metal3 s 0 50948 800 51188 6 la1_oenb[9]
port 211 nsew signal input
rlabel metal4 s 4208 2128 4528 57712 6 vccd1
port 212 nsew power input
rlabel metal4 s 34928 2128 35248 57712 6 vccd1
port 212 nsew power input
rlabel metal4 s 19568 2128 19888 57712 6 vssd1
port 213 nsew ground input
rlabel metal4 s 50288 2128 50608 57712 6 vssd1
port 213 nsew ground input
rlabel metal3 s 59200 27828 60000 28068 6 wb_clk_i
port 214 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 13677170
string GDS_FILE /openlane/designs/wrapped_wavelet_transform/runs/RUN_2022.06.06_03.17.52/results/finishing/wrapped_wavelet_transform.magic.gds
string GDS_START 1011494
<< end >>

