* NGSPICE file created from wrapped_wavelet_transform.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s50_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

.subckt wrapped_wavelet_transform active io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29]
+ io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32]
+ io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5]
+ io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1]
+ io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27]
+ io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34]
+ io_out[35] io_out[36] io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] la1_data_in[0] la1_data_in[10] la1_data_in[11] la1_data_in[12]
+ la1_data_in[13] la1_data_in[14] la1_data_in[15] la1_data_in[16] la1_data_in[17]
+ la1_data_in[18] la1_data_in[19] la1_data_in[1] la1_data_in[20] la1_data_in[21] la1_data_in[22]
+ la1_data_in[23] la1_data_in[24] la1_data_in[25] la1_data_in[26] la1_data_in[27]
+ la1_data_in[28] la1_data_in[29] la1_data_in[2] la1_data_in[30] la1_data_in[31] la1_data_in[3]
+ la1_data_in[4] la1_data_in[5] la1_data_in[6] la1_data_in[7] la1_data_in[8] la1_data_in[9]
+ la1_data_out[0] la1_data_out[10] la1_data_out[11] la1_data_out[12] la1_data_out[13]
+ la1_data_out[14] la1_data_out[15] la1_data_out[16] la1_data_out[17] la1_data_out[18]
+ la1_data_out[19] la1_data_out[1] la1_data_out[20] la1_data_out[21] la1_data_out[22]
+ la1_data_out[23] la1_data_out[24] la1_data_out[25] la1_data_out[26] la1_data_out[27]
+ la1_data_out[28] la1_data_out[29] la1_data_out[2] la1_data_out[30] la1_data_out[31]
+ la1_data_out[3] la1_data_out[4] la1_data_out[5] la1_data_out[6] la1_data_out[7]
+ la1_data_out[8] la1_data_out[9] la1_oenb[0] la1_oenb[10] la1_oenb[11] la1_oenb[12]
+ la1_oenb[13] la1_oenb[14] la1_oenb[15] la1_oenb[16] la1_oenb[17] la1_oenb[18] la1_oenb[19]
+ la1_oenb[1] la1_oenb[20] la1_oenb[21] la1_oenb[22] la1_oenb[23] la1_oenb[24] la1_oenb[25]
+ la1_oenb[26] la1_oenb[27] la1_oenb[28] la1_oenb[29] la1_oenb[2] la1_oenb[30] la1_oenb[31]
+ la1_oenb[3] la1_oenb[4] la1_oenb[5] la1_oenb[6] la1_oenb[7] la1_oenb[8] la1_oenb[9]
+ vccd1 vssd1 wb_clk_i
XFILLER_100_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6914_ hold61/A _6893_/B _6894_/A hold65/X vssd1 vssd1 vccd1 vccd1 _6914_/X sky130_fd_sc_hd__a22o_1
XFILLER_23_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6845_ _6845_/A hold68/X vssd1 vssd1 vccd1 vccd1 hold67/A sky130_fd_sc_hd__or2_1
X_3988_ _7193_/Q vssd1 vssd1 vccd1 vccd1 _4694_/A sky130_fd_sc_hd__buf_2
XFILLER_10_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6776_ _6809_/A _6809_/B vssd1 vssd1 vccd1 vccd1 _6777_/B sky130_fd_sc_hd__xor2_1
X_5727_ _5727_/A _5728_/B vssd1 vssd1 vccd1 vccd1 _5760_/B sky130_fd_sc_hd__xor2_2
XFILLER_50_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5658_ _6938_/A _6679_/B vssd1 vssd1 vccd1 vccd1 _5692_/A sky130_fd_sc_hd__xnor2_2
X_4609_ _4609_/A _4609_/B vssd1 vssd1 vccd1 vccd1 _4616_/A sky130_fd_sc_hd__xnor2_1
X_5589_ _5589_/A _5589_/B vssd1 vssd1 vccd1 vccd1 _5590_/B sky130_fd_sc_hd__xnor2_1
XFILLER_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7328_ _7328_/A _3739_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[2] sky130_fd_sc_hd__ebufn_8
XFILLER_89_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7263__56 vssd1 vssd1 vccd1 vccd1 _7263__56/HI _7362_/A sky130_fd_sc_hd__conb_1
XFILLER_36_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4960_ hold99/A _3818_/B _3816_/X vssd1 vssd1 vccd1 vccd1 _5286_/B sky130_fd_sc_hd__a21oi_2
XFILLER_17_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4891_ _4891_/A _4891_/B vssd1 vssd1 vccd1 vccd1 _4892_/B sky130_fd_sc_hd__or2_1
X_3911_ _4957_/A _3998_/B _3865_/X vssd1 vssd1 vccd1 vccd1 _3912_/B sky130_fd_sc_hd__a21oi_1
X_3842_ _7187_/Q _7186_/Q vssd1 vssd1 vccd1 vccd1 _4506_/A sky130_fd_sc_hd__or2_2
X_6630_ _6628_/A _6628_/B _6656_/A vssd1 vssd1 vccd1 vccd1 _6631_/B sky130_fd_sc_hd__o21ba_1
X_6561_ _6559_/X _6560_/X _6417_/Y vssd1 vssd1 vccd1 vccd1 _6584_/B sky130_fd_sc_hd__a21oi_4
X_5512_ _5513_/A _5513_/B _5513_/C vssd1 vssd1 vccd1 vccd1 _5558_/B sky130_fd_sc_hd__o21ai_1
X_3773_ _5347_/A _7183_/Q vssd1 vssd1 vccd1 vccd1 _4285_/A sky130_fd_sc_hd__and2_2
X_6492_ _6492_/A _6492_/B vssd1 vssd1 vccd1 vccd1 _6520_/A sky130_fd_sc_hd__xnor2_4
X_5443_ _5444_/A _5444_/B vssd1 vssd1 vccd1 vccd1 _5575_/A sky130_fd_sc_hd__nand2_2
XFILLER_99_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5374_ _5380_/A _5380_/B vssd1 vssd1 vccd1 vccd1 _5375_/C sky130_fd_sc_hd__xnor2_1
X_7113_ _5391_/B _6933_/B _7112_/X _6405_/X vssd1 vssd1 vccd1 vccd1 _7222_/D sky130_fd_sc_hd__o211a_1
X_4325_ _4465_/B _4325_/B vssd1 vssd1 vccd1 vccd1 _4436_/A sky130_fd_sc_hd__xnor2_4
X_4256_ _4257_/A _4257_/B vssd1 vssd1 vccd1 vccd1 _4497_/B sky130_fd_sc_hd__xnor2_2
X_7044_ hold121/X _7032_/X _7043_/X _7034_/X vssd1 vssd1 vccd1 vccd1 _7195_/D sky130_fd_sc_hd__o211a_1
X_4187_ _4187_/A _4187_/B vssd1 vssd1 vccd1 vccd1 _4188_/B sky130_fd_sc_hd__xnor2_2
XFILLER_55_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6828_ _6828_/A _6828_/B vssd1 vssd1 vccd1 vccd1 _6831_/A sky130_fd_sc_hd__xnor2_1
X_6759_ _6758_/B _6759_/B vssd1 vssd1 vccd1 vccd1 _6760_/B sky130_fd_sc_hd__and2b_1
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5090_ _5091_/A _5091_/B vssd1 vssd1 vccd1 vccd1 _5092_/A sky130_fd_sc_hd__nor2_1
X_4110_ _4110_/A _4138_/B vssd1 vssd1 vccd1 vccd1 _6713_/A sky130_fd_sc_hd__nor2_4
X_4041_ _4120_/A _4120_/B vssd1 vssd1 vccd1 vccd1 _4237_/A sky130_fd_sc_hd__xnor2_4
XFILLER_68_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5992_ _6577_/A vssd1 vssd1 vccd1 vccd1 _6971_/A sky130_fd_sc_hd__buf_2
X_4943_ _4935_/X _4938_/X _4939_/Y _4940_/X _4942_/A vssd1 vssd1 vccd1 vccd1 _5111_/B
+ sky130_fd_sc_hd__a311o_4
X_4874_ _5873_/A vssd1 vssd1 vccd1 vccd1 _7014_/A sky130_fd_sc_hd__buf_2
X_6613_ _6613_/A _6613_/B vssd1 vssd1 vccd1 vccd1 _6619_/A sky130_fd_sc_hd__xnor2_1
X_3825_ _3825_/A vssd1 vssd1 vccd1 vccd1 _4527_/A sky130_fd_sc_hd__buf_2
X_6544_ _6544_/A _6544_/B vssd1 vssd1 vccd1 vccd1 _6546_/B sky130_fd_sc_hd__xor2_2
X_3756_ _7171_/Q _4789_/B vssd1 vssd1 vccd1 vccd1 _3805_/A sky130_fd_sc_hd__nand2_1
XFILLER_20_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6475_ _6475_/A _6475_/B _6475_/C _6475_/D vssd1 vssd1 vccd1 vccd1 _6475_/X sky130_fd_sc_hd__and4_1
X_3687_ _3691_/A vssd1 vssd1 vccd1 vccd1 _3687_/Y sky130_fd_sc_hd__inv_2
X_5426_ _5428_/A _5426_/B vssd1 vssd1 vccd1 vccd1 _5895_/A sky130_fd_sc_hd__nand2_2
X_5357_ _5420_/A _5357_/B vssd1 vssd1 vccd1 vccd1 _5358_/B sky130_fd_sc_hd__xnor2_1
X_4308_ _5932_/A _4308_/B vssd1 vssd1 vccd1 vccd1 _4460_/A sky130_fd_sc_hd__nand2b_2
XFILLER_59_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5288_ _5289_/A _5289_/B _5289_/C vssd1 vssd1 vccd1 vccd1 _5290_/A sky130_fd_sc_hd__a21oi_1
XFILLER_101_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4239_ _4239_/A _4239_/B vssd1 vssd1 vccd1 vccd1 _4494_/A sky130_fd_sc_hd__and2_2
X_7027_ _7063_/A vssd1 vssd1 vccd1 vccd1 _7038_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7233__26 vssd1 vssd1 vccd1 vccd1 _7233__26/HI _7332_/A sky130_fd_sc_hd__conb_1
X_7312__105 vssd1 vssd1 vccd1 vccd1 _7312__105/HI _7420_/A sky130_fd_sc_hd__conb_1
XFILLER_64_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4590_ hold91/A _6624_/A vssd1 vssd1 vccd1 vccd1 _4838_/A sky130_fd_sc_hd__xor2_2
X_3610_ _3734_/A vssd1 vssd1 vccd1 vccd1 _3742_/A sky130_fd_sc_hd__buf_4
X_6260_ _5594_/X hold114/X _5595_/X _6259_/X vssd1 vssd1 vccd1 vccd1 _7131_/D sky130_fd_sc_hd__o211a_1
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5211_ _5210_/A _5210_/B hold84/A vssd1 vssd1 vccd1 vccd1 _5335_/B sky130_fd_sc_hd__o21a_1
X_6191_ _6255_/A _6191_/B vssd1 vssd1 vccd1 vccd1 _6194_/A sky130_fd_sc_hd__xor2_4
XFILLER_69_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5142_ _5142_/A _5142_/B vssd1 vssd1 vccd1 vccd1 _5151_/A sky130_fd_sc_hd__nand2_1
XFILLER_96_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5073_ _5339_/A _5073_/B vssd1 vssd1 vccd1 vccd1 _5073_/Y sky130_fd_sc_hd__nor2_1
X_4024_ _4024_/A _4024_/B vssd1 vssd1 vccd1 vccd1 _4025_/B sky130_fd_sc_hd__xnor2_2
XFILLER_37_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5975_ _5975_/A _5975_/B vssd1 vssd1 vccd1 vccd1 _5999_/B sky130_fd_sc_hd__xor2_1
X_4926_ _4888_/A _4888_/B _4925_/X vssd1 vssd1 vccd1 vccd1 _4926_/Y sky130_fd_sc_hd__a21oi_1
X_4857_ hold80/A _4857_/B vssd1 vssd1 vccd1 vccd1 _4895_/A sky130_fd_sc_hd__nand2_2
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3808_ _4481_/A _4481_/B vssd1 vssd1 vccd1 vccd1 _4485_/A sky130_fd_sc_hd__nor2_1
X_4788_ _4788_/A _4788_/B vssd1 vssd1 vccd1 vccd1 _4837_/A sky130_fd_sc_hd__xnor2_1
X_6527_ _6852_/A _6527_/B vssd1 vssd1 vccd1 vccd1 _6737_/A sky130_fd_sc_hd__xnor2_1
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3739_ _3739_/A vssd1 vssd1 vccd1 vccd1 _3739_/Y sky130_fd_sc_hd__inv_2
X_6458_ _6458_/A _6458_/B _6727_/A vssd1 vssd1 vccd1 vccd1 _6459_/B sky130_fd_sc_hd__and3_1
X_6389_ _6359_/A _6359_/B _6388_/X vssd1 vssd1 vccd1 vccd1 _6390_/B sky130_fd_sc_hd__a21o_1
X_5409_ _6524_/A _5409_/B vssd1 vssd1 vccd1 vccd1 _5412_/C sky130_fd_sc_hd__nand2_1
X_7299__92 vssd1 vssd1 vccd1 vccd1 _7299__92/HI _7407_/A sky130_fd_sc_hd__conb_1
XFILLER_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5760_ _5760_/A _5760_/B vssd1 vssd1 vccd1 vccd1 _5774_/A sky130_fd_sc_hd__xor2_2
XFILLER_22_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4711_ _4710_/A _4711_/B vssd1 vssd1 vccd1 vccd1 _4711_/X sky130_fd_sc_hd__and2b_1
X_5691_ _6484_/B _5691_/B vssd1 vssd1 vccd1 vccd1 _5721_/A sky130_fd_sc_hd__nand2_2
X_7430_ _7430_/A _3729_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[34] sky130_fd_sc_hd__ebufn_8
X_4642_ _4642_/A _4642_/B vssd1 vssd1 vccd1 vccd1 _4650_/B sky130_fd_sc_hd__xnor2_1
X_7361_ _7361_/A _3625_/Y vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__ebufn_8
X_4573_ _4573_/A _4795_/B vssd1 vssd1 vccd1 vccd1 _5850_/B sky130_fd_sc_hd__nor2_1
X_6312_ _6828_/A _6243_/B _6244_/A _6311_/X vssd1 vssd1 vccd1 vccd1 _6313_/B sky130_fd_sc_hd__a31o_1
X_6243_ _6413_/A _6243_/B vssd1 vssd1 vccd1 vccd1 _6244_/B sky130_fd_sc_hd__nand2_1
X_6174_ _6174_/A vssd1 vssd1 vccd1 vccd1 _6962_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_97_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5125_ _5125_/A _5267_/B vssd1 vssd1 vccd1 vccd1 _5127_/C sky130_fd_sc_hd__xnor2_1
XFILLER_57_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5056_ hold58/A _5056_/B _5056_/C _5056_/D vssd1 vssd1 vccd1 vccd1 _5067_/B sky130_fd_sc_hd__or4_1
X_4007_ _4007_/A _4007_/B vssd1 vssd1 vccd1 vccd1 _4240_/B sky130_fd_sc_hd__xnor2_1
XFILLER_72_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5958_ _5963_/A _5963_/B vssd1 vssd1 vccd1 vccd1 _5965_/A sky130_fd_sc_hd__and2b_1
XFILLER_13_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4909_ _5644_/A _6678_/A vssd1 vssd1 vccd1 vccd1 _4910_/B sky130_fd_sc_hd__or2_1
XFILLER_40_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5889_ _5890_/A _5890_/B vssd1 vssd1 vccd1 vccd1 _5894_/B sky130_fd_sc_hd__xor2_1
XFILLER_20_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__clkbuf_2
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_75_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold85 hold85/A vssd1 vssd1 vccd1 vccd1 hold85/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_28_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_5 _5165_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7318__111 vssd1 vssd1 vccd1 vccd1 _7318__111/HI _7426_/A sky130_fd_sc_hd__conb_1
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6930_ input2/X _7116_/B _6929_/Y _6846_/X vssd1 vssd1 vccd1 vccd1 _7153_/D sky130_fd_sc_hd__o211a_1
XFILLER_81_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6861_ _6862_/A _6862_/B _6862_/C vssd1 vssd1 vccd1 vccd1 _6875_/B sky130_fd_sc_hd__o21ai_1
XFILLER_34_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5812_ _5812_/A _5812_/B vssd1 vssd1 vccd1 vccd1 _5813_/B sky130_fd_sc_hd__xnor2_1
X_6792_ _6792_/A _6792_/B vssd1 vssd1 vccd1 vccd1 _6814_/A sky130_fd_sc_hd__or2_1
XFILLER_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5743_ _6054_/A _5743_/B vssd1 vssd1 vccd1 vccd1 _5744_/B sky130_fd_sc_hd__nand2_1
X_5674_ _7190_/Q _5674_/B vssd1 vssd1 vccd1 vccd1 _5676_/A sky130_fd_sc_hd__and2b_1
X_4625_ _4625_/A _4626_/B vssd1 vssd1 vccd1 vccd1 _4688_/B sky130_fd_sc_hd__xnor2_1
X_7413_ _7413_/A _3733_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[17] sky130_fd_sc_hd__ebufn_8
X_7344_ _7344_/A _3628_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[18] sky130_fd_sc_hd__ebufn_8
X_4556_ _4556_/A _4556_/B vssd1 vssd1 vccd1 vccd1 _4652_/B sky130_fd_sc_hd__or2_1
XFILLER_89_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4487_ _6120_/A _4487_/B vssd1 vssd1 vccd1 vccd1 _4562_/B sky130_fd_sc_hd__xor2_4
X_6226_ _6575_/A _6226_/B vssd1 vssd1 vccd1 vccd1 _6302_/A sky130_fd_sc_hd__nand2_1
X_7269__62 vssd1 vssd1 vccd1 vccd1 _7269__62/HI _7368_/A sky130_fd_sc_hd__conb_1
XFILLER_85_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6157_ _6539_/A vssd1 vssd1 vccd1 vccd1 _6528_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5108_ _5108_/A _5108_/B vssd1 vssd1 vccd1 vccd1 _5108_/X sky130_fd_sc_hd__and2_1
XFILLER_85_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6088_ _6088_/A _6088_/B vssd1 vssd1 vccd1 vccd1 _6089_/B sky130_fd_sc_hd__nor2_2
X_5039_ _5039_/A _4045_/A vssd1 vssd1 vccd1 vccd1 _5039_/X sky130_fd_sc_hd__or2b_1
XFILLER_26_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4410_ _4412_/A _4799_/A vssd1 vssd1 vccd1 vccd1 _4649_/B sky130_fd_sc_hd__nand2_1
X_5390_ _5391_/A _5391_/B _5287_/A vssd1 vssd1 vccd1 vccd1 _5541_/B sky130_fd_sc_hd__a21oi_2
XFILLER_99_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4341_ _4338_/A _4338_/B _4443_/A vssd1 vssd1 vccd1 vccd1 _5101_/B sky130_fd_sc_hd__o21ai_4
X_7060_ _7073_/A vssd1 vssd1 vccd1 vccd1 _7060_/X sky130_fd_sc_hd__clkbuf_2
X_4272_ _4272_/A _5707_/B vssd1 vssd1 vccd1 vccd1 _4272_/X sky130_fd_sc_hd__or2_1
X_6011_ _6011_/A _6011_/B vssd1 vssd1 vccd1 vccd1 _6011_/Y sky130_fd_sc_hd__nand2_1
XFILLER_94_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6913_ _7116_/A hold4/X vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__nor2_1
XFILLER_23_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6844_ _6844_/A _6869_/B vssd1 vssd1 vccd1 vccd1 _6844_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3987_ _4638_/B _3993_/B vssd1 vssd1 vccd1 vccd1 _4014_/A sky130_fd_sc_hd__xnor2_2
XFILLER_22_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6775_ _6740_/A _6740_/B _6774_/X vssd1 vssd1 vccd1 vccd1 _6809_/B sky130_fd_sc_hd__a21bo_1
X_5726_ _5762_/A _5762_/B _5725_/X vssd1 vssd1 vccd1 vccd1 _5728_/B sky130_fd_sc_hd__a21bo_1
X_5657_ _6483_/B vssd1 vssd1 vccd1 vccd1 _6466_/A sky130_fd_sc_hd__clkbuf_2
X_4608_ _4608_/A _4608_/B vssd1 vssd1 vccd1 vccd1 _4700_/A sky130_fd_sc_hd__xor2_1
X_5588_ _5588_/A _5588_/B vssd1 vssd1 vccd1 vccd1 _5589_/B sky130_fd_sc_hd__xnor2_1
X_4539_ _4539_/A _4539_/B _4539_/C vssd1 vssd1 vccd1 vccd1 _4539_/X sky130_fd_sc_hd__or3_1
X_7327_ _7327_/A _3738_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[1] sky130_fd_sc_hd__ebufn_8
XFILLER_7_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6209_ _6209_/A _6264_/B vssd1 vssd1 vccd1 vccd1 _6212_/A sky130_fd_sc_hd__xnor2_2
X_7189_ _7222_/CLK _7189_/D vssd1 vssd1 vccd1 vccd1 _7189_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4890_ _4890_/A _4890_/B vssd1 vssd1 vccd1 vccd1 _4904_/A sky130_fd_sc_hd__or2_1
XFILLER_83_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3910_ _3910_/A _3998_/B vssd1 vssd1 vccd1 vccd1 _3912_/A sky130_fd_sc_hd__xnor2_1
X_3841_ _4613_/A _4249_/A vssd1 vssd1 vccd1 vccd1 _4011_/B sky130_fd_sc_hd__nor2_1
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3772_ _7190_/Q vssd1 vssd1 vccd1 vccd1 _5347_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6560_ _6560_/A _6411_/B vssd1 vssd1 vccd1 vccd1 _6560_/X sky130_fd_sc_hd__or2b_1
X_5511_ _5558_/A _5511_/B vssd1 vssd1 vccd1 vccd1 _5513_/C sky130_fd_sc_hd__and2_1
X_6491_ _6491_/A _6491_/B vssd1 vssd1 vccd1 vccd1 _6492_/A sky130_fd_sc_hd__nand2_2
X_5442_ _5442_/A _5442_/B vssd1 vssd1 vccd1 vccd1 _5444_/B sky130_fd_sc_hd__nor2_1
X_5373_ _5253_/A _5253_/B _5372_/Y vssd1 vssd1 vccd1 vccd1 _5380_/B sky130_fd_sc_hd__o21a_1
X_4324_ _4316_/A _4316_/B _4323_/X vssd1 vssd1 vccd1 vccd1 _4445_/A sky130_fd_sc_hd__o21ai_4
X_7112_ hold96/X _7114_/B vssd1 vssd1 vccd1 vccd1 _7112_/X sky130_fd_sc_hd__or2_1
XFILLER_87_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7043_ _7043_/A _7059_/B vssd1 vssd1 vccd1 vccd1 _7043_/X sky130_fd_sc_hd__or2_1
X_7239__32 vssd1 vssd1 vccd1 vccd1 _7239__32/HI _7338_/A sky130_fd_sc_hd__conb_1
X_4255_ _4500_/A _4500_/B _4254_/X vssd1 vssd1 vccd1 vccd1 _4257_/B sky130_fd_sc_hd__a21oi_1
XFILLER_86_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4186_ _4243_/A _4243_/B _4185_/X vssd1 vssd1 vccd1 vccd1 _4188_/A sky130_fd_sc_hd__a21oi_2
XFILLER_94_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6827_ _6827_/A _6827_/B vssd1 vssd1 vccd1 vccd1 _6828_/B sky130_fd_sc_hd__xnor2_1
XFILLER_23_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6758_ _6759_/B _6758_/B vssd1 vssd1 vccd1 vccd1 _6812_/A sky130_fd_sc_hd__and2b_1
X_6689_ _6947_/A _6693_/B vssd1 vssd1 vccd1 vccd1 _6690_/B sky130_fd_sc_hd__or2_1
X_5709_ _5709_/A _5709_/B vssd1 vssd1 vccd1 vccd1 _5710_/B sky130_fd_sc_hd__nor2_2
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4040_ _4187_/A _4187_/B _4039_/X vssd1 vssd1 vccd1 vccd1 _4120_/B sky130_fd_sc_hd__a21oi_2
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5991_ _5991_/A vssd1 vssd1 vccd1 vccd1 _6950_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_64_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4942_ _4942_/A _4942_/B vssd1 vssd1 vccd1 vccd1 _4942_/Y sky130_fd_sc_hd__nand2_2
X_4873_ _4873_/A vssd1 vssd1 vccd1 vccd1 _5873_/A sky130_fd_sc_hd__buf_2
XFILLER_60_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6612_ _6711_/A _6711_/B vssd1 vssd1 vccd1 vccd1 _6647_/A sky130_fd_sc_hd__xnor2_2
X_3824_ _5129_/A vssd1 vssd1 vccd1 vccd1 _5273_/A sky130_fd_sc_hd__inv_2
XFILLER_20_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6543_ _6480_/A _6480_/B _6480_/C _6565_/B _6510_/X vssd1 vssd1 vccd1 vccd1 _6544_/B
+ sky130_fd_sc_hd__a41o_1
X_3755_ _7168_/Q vssd1 vssd1 vccd1 vccd1 _4789_/B sky130_fd_sc_hd__clkbuf_2
X_6474_ _6725_/A _6725_/B vssd1 vssd1 vccd1 vccd1 _6765_/B sky130_fd_sc_hd__nand2_1
X_3686_ _3710_/A vssd1 vssd1 vccd1 vccd1 _3691_/A sky130_fd_sc_hd__buf_12
X_5425_ _6564_/A _5737_/A vssd1 vssd1 vccd1 vccd1 _5426_/B sky130_fd_sc_hd__or2_1
XFILLER_99_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5356_ _5356_/A _5356_/B vssd1 vssd1 vccd1 vccd1 _5357_/B sky130_fd_sc_hd__xor2_1
XFILLER_101_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4307_ _4329_/A _4795_/A vssd1 vssd1 vccd1 vccd1 _4308_/B sky130_fd_sc_hd__nand2_1
XFILLER_59_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5287_ _5287_/A _5287_/B vssd1 vssd1 vccd1 vccd1 _5289_/C sky130_fd_sc_hd__xnor2_1
X_4238_ _4238_/A _4238_/B vssd1 vssd1 vccd1 vccd1 _4239_/B sky130_fd_sc_hd__nand2_1
X_7026_ _7003_/A _7018_/X _7025_/X _7021_/X vssd1 vssd1 vccd1 vccd1 _7188_/D sky130_fd_sc_hd__o211a_1
XFILLER_28_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4169_ _4799_/B vssd1 vssd1 vccd1 vccd1 _4857_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_74_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5210_ _5210_/A _5210_/B vssd1 vssd1 vccd1 vccd1 _5210_/Y sky130_fd_sc_hd__nand2_1
X_6190_ _6096_/A _6096_/B _6189_/X vssd1 vssd1 vccd1 vccd1 _6191_/B sky130_fd_sc_hd__o21ai_4
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5141_ _5141_/A _5141_/B _5141_/C vssd1 vssd1 vccd1 vccd1 _5142_/B sky130_fd_sc_hd__or3_1
X_5072_ _5218_/A vssd1 vssd1 vccd1 vccd1 _5339_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4023_ _4021_/X _4007_/B _4022_/X vssd1 vssd1 vccd1 vccd1 _4025_/A sky130_fd_sc_hd__o21a_1
XFILLER_77_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5974_ _5953_/B _5973_/X _5596_/A vssd1 vssd1 vccd1 vccd1 _5981_/B sky130_fd_sc_hd__a21bo_1
XFILLER_40_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4925_ _4887_/B _4925_/B vssd1 vssd1 vccd1 vccd1 _4925_/X sky130_fd_sc_hd__and2b_1
X_4856_ _4856_/A _4856_/B vssd1 vssd1 vccd1 vccd1 _4858_/B sky130_fd_sc_hd__nor2_1
X_3807_ _3807_/A _3807_/B vssd1 vssd1 vccd1 vccd1 _4481_/B sky130_fd_sc_hd__nor2_1
X_4787_ _4787_/A _4787_/B vssd1 vssd1 vccd1 vccd1 _4787_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_20_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6526_ _6526_/A _6733_/B vssd1 vssd1 vccd1 vccd1 _6527_/B sky130_fd_sc_hd__xnor2_2
X_3738_ _3739_/A vssd1 vssd1 vccd1 vccd1 _3738_/Y sky130_fd_sc_hd__inv_2
X_3669_ _3672_/A vssd1 vssd1 vccd1 vccd1 _3669_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6457_ _6727_/A _6457_/B vssd1 vssd1 vccd1 vccd1 _6728_/A sky130_fd_sc_hd__and2b_1
X_6388_ _6356_/A _6388_/B vssd1 vssd1 vccd1 vccd1 _6388_/X sky130_fd_sc_hd__and2b_1
X_5408_ _6523_/A vssd1 vssd1 vccd1 vccd1 _6524_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_87_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5339_ _5339_/A _5339_/B vssd1 vssd1 vccd1 vccd1 _5446_/C sky130_fd_sc_hd__xor2_1
XFILLER_85_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7009_ _7009_/A _7011_/B vssd1 vssd1 vccd1 vccd1 _7009_/X sky130_fd_sc_hd__or2_1
XFILLER_90_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4710_ _4710_/A _4711_/B vssd1 vssd1 vccd1 vccd1 _4756_/B sky130_fd_sc_hd__xnor2_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5690_ _5690_/A _7175_/Q vssd1 vssd1 vccd1 vccd1 _5715_/B sky130_fd_sc_hd__or2_1
X_4641_ _4641_/A _4641_/B vssd1 vssd1 vccd1 vccd1 _4642_/B sky130_fd_sc_hd__nor2_1
X_4572_ _4572_/A _4795_/B vssd1 vssd1 vccd1 vccd1 _4744_/B sky130_fd_sc_hd__and2_1
X_7360_ _7360_/A _3635_/Y vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__ebufn_8
X_6311_ _6245_/A _6311_/B vssd1 vssd1 vccd1 vccd1 _6311_/X sky130_fd_sc_hd__and2b_1
X_6242_ _6301_/A _6960_/A vssd1 vssd1 vccd1 vccd1 _6243_/B sky130_fd_sc_hd__or2b_1
X_6173_ _6173_/A _6247_/A vssd1 vssd1 vccd1 vccd1 _6182_/A sky130_fd_sc_hd__xnor2_4
XFILLER_97_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5124_ _5124_/A _5394_/A vssd1 vssd1 vccd1 vccd1 _5267_/B sky130_fd_sc_hd__and2_1
XFILLER_57_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5055_ _5055_/A _5056_/D vssd1 vssd1 vccd1 vccd1 _5067_/A sky130_fd_sc_hd__or2_1
X_4006_ _4002_/A _4002_/B _4005_/X vssd1 vssd1 vccd1 vccd1 _4007_/B sky130_fd_sc_hd__o21a_1
XFILLER_65_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5957_ _5957_/A _6002_/A vssd1 vssd1 vccd1 vccd1 _5963_/B sky130_fd_sc_hd__nand2_1
X_4908_ _5880_/B vssd1 vssd1 vccd1 vccd1 _5987_/A sky130_fd_sc_hd__buf_2
X_5888_ _5907_/A _5907_/B _5887_/A vssd1 vssd1 vccd1 vccd1 _5890_/B sky130_fd_sc_hd__a21oi_2
XFILLER_21_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4839_ _4838_/A _4838_/B _4838_/C vssd1 vssd1 vccd1 vccd1 _4839_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_21_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6509_ _6505_/A _6505_/B _6505_/C vssd1 vssd1 vccd1 vccd1 _6542_/B sky130_fd_sc_hd__a21o_1
XFILLER_20_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold64 hold64/A vssd1 vssd1 vccd1 vccd1 hold64/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold86/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold75 hold75/A vssd1 vssd1 vccd1 vccd1 hold75/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_90_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_6 _5200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6860_ _6875_/A _6860_/B vssd1 vssd1 vccd1 vccd1 _6862_/C sky130_fd_sc_hd__and2_1
XFILLER_34_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6791_ _5594_/X hold17/X _5595_/X _6790_/X vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__o211a_1
X_5811_ _5811_/A _5811_/B vssd1 vssd1 vccd1 vccd1 _6092_/A sky130_fd_sc_hd__xnor2_2
X_5742_ _6620_/A _5756_/A vssd1 vssd1 vccd1 vccd1 _5743_/B sky130_fd_sc_hd__nand2_1
X_5673_ _5673_/A _5673_/B _5673_/C vssd1 vssd1 vccd1 vccd1 _5685_/A sky130_fd_sc_hd__and3_1
X_4624_ _4690_/A _4690_/B _4623_/X vssd1 vssd1 vccd1 vccd1 _4626_/B sky130_fd_sc_hd__a21bo_1
X_7412_ _7412_/A _3708_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[16] sky130_fd_sc_hd__ebufn_8
X_4555_ _4555_/A _4555_/B vssd1 vssd1 vccd1 vccd1 _4556_/B sky130_fd_sc_hd__and2_1
X_7343_ _7343_/A _3627_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[17] sky130_fd_sc_hd__ebufn_8
X_4486_ _4486_/A _4486_/B vssd1 vssd1 vccd1 vccd1 _4487_/B sky130_fd_sc_hd__xnor2_2
X_6225_ _6298_/A _6298_/B vssd1 vssd1 vccd1 vccd1 _6235_/A sky130_fd_sc_hd__xor2_4
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6156_ _6156_/A _6236_/B vssd1 vssd1 vccd1 vccd1 _6170_/A sky130_fd_sc_hd__xor2_4
XFILLER_85_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5107_ _5107_/A _5107_/B vssd1 vssd1 vccd1 vccd1 _5110_/A sky130_fd_sc_hd__xnor2_2
X_7284__77 vssd1 vssd1 vccd1 vccd1 _7284__77/HI _7392_/A sky130_fd_sc_hd__conb_1
XFILLER_85_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6087_ _6805_/A _6087_/B vssd1 vssd1 vccd1 vccd1 _6088_/B sky130_fd_sc_hd__nor2_1
X_5038_ _5183_/A _5183_/B vssd1 vssd1 vccd1 vccd1 _5243_/A sky130_fd_sc_hd__xnor2_1
XFILLER_45_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6989_ _7063_/A vssd1 vssd1 vccd1 vccd1 _7011_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_25_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4340_ _4442_/A _4442_/B vssd1 vssd1 vccd1 vccd1 _4443_/A sky130_fd_sc_hd__nand2_1
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4271_ _4272_/A _5707_/B vssd1 vssd1 vccd1 vccd1 _4315_/B sky130_fd_sc_hd__xnor2_2
XFILLER_79_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6010_ _6011_/A _6011_/B vssd1 vssd1 vccd1 vccd1 _6010_/X sky130_fd_sc_hd__or2_1
XFILLER_39_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6912_ hold2/X _6893_/A _6911_/X vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__a21oi_1
X_6843_ _6786_/A _6789_/Y _6840_/Y _6816_/B _6842_/A vssd1 vssd1 vccd1 vccd1 _6869_/B
+ sky130_fd_sc_hd__a311oi_2
XFILLER_35_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3986_ _4533_/A _3986_/B vssd1 vssd1 vccd1 vccd1 _3993_/B sky130_fd_sc_hd__xnor2_2
X_6774_ _6774_/A _6739_/A vssd1 vssd1 vccd1 vccd1 _6774_/X sky130_fd_sc_hd__or2b_1
X_5725_ _5725_/A _5724_/B vssd1 vssd1 vccd1 vccd1 _5725_/X sky130_fd_sc_hd__or2b_1
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5656_ _6014_/A _6014_/B vssd1 vssd1 vccd1 vccd1 _5682_/A sky130_fd_sc_hd__xor2_2
X_4607_ _4607_/A _4607_/B vssd1 vssd1 vccd1 vccd1 _4619_/A sky130_fd_sc_hd__xnor2_2
X_5587_ _5587_/A _5587_/B vssd1 vssd1 vccd1 vccd1 _5588_/B sky130_fd_sc_hd__xnor2_1
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4538_ _4538_/A _4538_/B vssd1 vssd1 vccd1 vccd1 _4539_/C sky130_fd_sc_hd__xor2_1
X_7326_ _7326_/A _3737_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[0] sky130_fd_sc_hd__ebufn_8
XFILLER_2_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4469_ _6410_/A _4469_/B _4469_/C vssd1 vssd1 vccd1 vccd1 _4566_/A sky130_fd_sc_hd__and3_1
X_6208_ _6263_/A _6263_/B vssd1 vssd1 vccd1 vccd1 _6264_/B sky130_fd_sc_hd__xor2_2
X_7188_ _7221_/CLK _7188_/D vssd1 vssd1 vccd1 vccd1 _7188_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_58_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6139_ _6139_/A vssd1 vssd1 vccd1 vccd1 _6329_/A sky130_fd_sc_hd__clkbuf_2
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3840_ _7188_/Q _5674_/B vssd1 vssd1 vccd1 vccd1 _4249_/A sky130_fd_sc_hd__xor2_2
XFILLER_32_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3771_ _3801_/A _3801_/B _3770_/Y vssd1 vssd1 vccd1 vccd1 _3798_/A sky130_fd_sc_hd__o21ai_2
X_5510_ _5510_/A _5510_/B _5510_/C vssd1 vssd1 vccd1 vccd1 _5511_/B sky130_fd_sc_hd__or3_1
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6490_ _6514_/A _6514_/B vssd1 vssd1 vccd1 vccd1 _6490_/X sky130_fd_sc_hd__and2_1
X_5441_ _5547_/A _5547_/B vssd1 vssd1 vccd1 vccd1 _5442_/B sky130_fd_sc_hd__and2_1
XFILLER_99_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5372_ _5372_/A _5372_/B vssd1 vssd1 vccd1 vccd1 _5372_/Y sky130_fd_sc_hd__nand2_1
XFILLER_99_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4323_ _4456_/B _4456_/A vssd1 vssd1 vccd1 vccd1 _4323_/X sky130_fd_sc_hd__or2b_1
X_7111_ _7091_/A _7101_/X _7110_/X _6405_/X vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__o211a_1
X_7042_ _7019_/A _7032_/X _7041_/X _7034_/X vssd1 vssd1 vccd1 vccd1 _7194_/D sky130_fd_sc_hd__o211a_1
XFILLER_101_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4254_ _4253_/A _4254_/B vssd1 vssd1 vccd1 vccd1 _4254_/X sky130_fd_sc_hd__and2b_1
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4185_ _4185_/A _4185_/B vssd1 vssd1 vccd1 vccd1 _4185_/X sky130_fd_sc_hd__and2_1
XFILLER_86_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7254__47 vssd1 vssd1 vccd1 vccd1 _7254__47/HI _7353_/A sky130_fd_sc_hd__conb_1
XFILLER_55_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6826_ _6856_/A _6856_/B vssd1 vssd1 vccd1 vccd1 _6827_/B sky130_fd_sc_hd__or2_1
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6757_ _6720_/A _6720_/B _6723_/B vssd1 vssd1 vccd1 vccd1 _6759_/B sky130_fd_sc_hd__a21oi_1
XFILLER_23_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3969_ _6445_/B _7223_/Q vssd1 vssd1 vccd1 vccd1 _5023_/A sky130_fd_sc_hd__and2b_1
X_5708_ _5707_/B _5708_/B vssd1 vssd1 vccd1 vccd1 _5709_/B sky130_fd_sc_hd__and2b_1
X_6688_ _6688_/A _6688_/B vssd1 vssd1 vccd1 vccd1 _6693_/B sky130_fd_sc_hd__xnor2_1
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5639_ _5866_/A _5900_/A vssd1 vssd1 vccd1 vccd1 _5867_/A sky130_fd_sc_hd__nand2_1
XFILLER_2_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5990_ _5990_/A _5990_/B vssd1 vssd1 vccd1 vccd1 _5990_/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4941_ _4935_/X _4938_/X _4939_/Y _4940_/X vssd1 vssd1 vccd1 vccd1 _4942_/B sky130_fd_sc_hd__a31o_1
X_4872_ _4872_/A _4872_/B vssd1 vssd1 vccd1 vccd1 _4876_/A sky130_fd_sc_hd__nand2_1
X_3823_ _4956_/B vssd1 vssd1 vccd1 vccd1 _5129_/A sky130_fd_sc_hd__clkbuf_2
X_6611_ _6611_/A _6710_/A vssd1 vssd1 vccd1 vccd1 _6711_/B sky130_fd_sc_hd__xnor2_1
X_6542_ _6506_/C _6542_/B vssd1 vssd1 vccd1 vccd1 _6565_/B sky130_fd_sc_hd__and2b_1
X_3754_ _3754_/A vssd1 vssd1 vccd1 vccd1 _3770_/A sky130_fd_sc_hd__clkbuf_4
X_6473_ _6473_/A _6473_/B vssd1 vssd1 vccd1 vccd1 _6725_/B sky130_fd_sc_hd__xnor2_1
X_3685_ input1/X vssd1 vssd1 vccd1 vccd1 _3710_/A sky130_fd_sc_hd__clkbuf_4
X_5424_ _6564_/A _5737_/A vssd1 vssd1 vccd1 vccd1 _5428_/A sky130_fd_sc_hd__nand2_1
XFILLER_99_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5355_ _5355_/A _5355_/B vssd1 vssd1 vccd1 vccd1 _5356_/B sky130_fd_sc_hd__nor2_1
XFILLER_99_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4306_ _7163_/Q _7162_/Q _7161_/Q vssd1 vssd1 vccd1 vccd1 _5932_/A sky130_fd_sc_hd__o21a_1
XFILLER_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5286_ _5286_/A _5286_/B _5286_/C vssd1 vssd1 vccd1 vccd1 _5289_/A sky130_fd_sc_hd__or3_1
X_7025_ _7025_/A _7025_/B vssd1 vssd1 vccd1 vccd1 _7025_/X sky130_fd_sc_hd__or2_1
X_4237_ _4237_/A _4237_/B vssd1 vssd1 vccd1 vccd1 _4262_/A sky130_fd_sc_hd__xor2_4
XFILLER_67_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4168_ _7208_/Q vssd1 vssd1 vccd1 vccd1 _4799_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_83_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4099_ _7162_/Q _7161_/Q vssd1 vssd1 vccd1 vccd1 _4450_/B sky130_fd_sc_hd__xor2_4
XFILLER_28_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6809_ _6809_/A _6809_/B vssd1 vssd1 vccd1 vccd1 _6809_/Y sky130_fd_sc_hd__nand2_1
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5140_ _5141_/A _5141_/B _5141_/C vssd1 vssd1 vccd1 vccd1 _5142_/A sky130_fd_sc_hd__o21ai_1
XFILLER_96_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5071_ _5071_/A _5071_/B vssd1 vssd1 vccd1 vccd1 _5075_/A sky130_fd_sc_hd__xnor2_1
X_4022_ _4022_/A _3997_/B vssd1 vssd1 vccd1 vccd1 _4022_/X sky130_fd_sc_hd__or2b_1
XFILLER_49_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5973_ _6794_/A _6409_/B vssd1 vssd1 vccd1 vccd1 _5973_/X sky130_fd_sc_hd__or2_1
X_4924_ _4903_/A _4907_/X _4922_/X _4923_/X vssd1 vssd1 vccd1 vccd1 _4924_/X sky130_fd_sc_hd__o211a_1
XFILLER_52_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4855_ _4856_/A _4856_/B vssd1 vssd1 vccd1 vccd1 _4858_/A sky130_fd_sc_hd__and2_1
XFILLER_60_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4786_ _4786_/A vssd1 vssd1 vccd1 vccd1 _4787_/B sky130_fd_sc_hd__inv_2
X_3806_ _7066_/A hold98/A vssd1 vssd1 vccd1 vccd1 _3807_/B sky130_fd_sc_hd__nor2_1
X_3737_ _3739_/A vssd1 vssd1 vccd1 vccd1 _3737_/Y sky130_fd_sc_hd__inv_2
X_6525_ _6531_/A _6531_/B _6524_/X vssd1 vssd1 vccd1 vccd1 _6733_/B sky130_fd_sc_hd__a21o_1
X_3668_ _3672_/A vssd1 vssd1 vccd1 vccd1 _3668_/Y sky130_fd_sc_hd__inv_2
X_6456_ _6458_/A _6458_/B vssd1 vssd1 vccd1 vccd1 _6457_/B sky130_fd_sc_hd__nand2_1
X_6387_ _6393_/B _6387_/B vssd1 vssd1 vccd1 vccd1 _6390_/A sky130_fd_sc_hd__xnor2_1
X_5407_ _6523_/A _5409_/B vssd1 vssd1 vccd1 vccd1 _5412_/B sky130_fd_sc_hd__or2_1
X_5338_ _5423_/A _5423_/B vssd1 vssd1 vccd1 vccd1 _5339_/B sky130_fd_sc_hd__xnor2_1
XFILLER_87_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7008_ _6528_/B _7005_/X _7006_/Y _7007_/X vssd1 vssd1 vccd1 vccd1 _7181_/D sky130_fd_sc_hd__o211a_1
X_5269_ _5391_/A _5478_/A vssd1 vssd1 vccd1 vccd1 _5271_/B sky130_fd_sc_hd__xnor2_1
XFILLER_75_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4640_ _4695_/A _4695_/B vssd1 vssd1 vccd1 vccd1 _4650_/A sky130_fd_sc_hd__nor2_1
X_4571_ _7176_/Q vssd1 vssd1 vccd1 vccd1 _4914_/B sky130_fd_sc_hd__clkbuf_2
X_6310_ _6413_/A vssd1 vssd1 vccd1 vccd1 _6828_/A sky130_fd_sc_hd__buf_2
X_6241_ _6241_/A vssd1 vssd1 vccd1 vccd1 _6960_/A sky130_fd_sc_hd__buf_2
X_6172_ _6079_/A _6078_/A _6078_/B _6171_/X vssd1 vssd1 vccd1 vccd1 _6247_/A sky130_fd_sc_hd__o31a_2
XFILLER_97_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5123_ _5122_/B _5277_/B _5133_/A vssd1 vssd1 vccd1 vccd1 _5394_/A sky130_fd_sc_hd__o21ai_2
XFILLER_57_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5054_ _5054_/A _5054_/B vssd1 vssd1 vccd1 vccd1 _5341_/A sky130_fd_sc_hd__xor2_4
X_4005_ _4176_/A _4176_/B vssd1 vssd1 vccd1 vccd1 _4005_/X sky130_fd_sc_hd__or2b_1
XFILLER_53_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5956_ _6001_/A _6001_/B vssd1 vssd1 vccd1 vccd1 _6002_/A sky130_fd_sc_hd__nand2_1
X_4907_ _4907_/A _4923_/A vssd1 vssd1 vccd1 vccd1 _4907_/X sky130_fd_sc_hd__xor2_1
X_5887_ _5887_/A _5887_/B vssd1 vssd1 vccd1 vccd1 _5907_/B sky130_fd_sc_hd__nor2_1
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4838_ _4838_/A _4838_/B _4838_/C vssd1 vssd1 vccd1 vccd1 _4838_/X sky130_fd_sc_hd__and3_1
XFILLER_21_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4769_ _4820_/A _4820_/B _4768_/X vssd1 vssd1 vccd1 vccd1 _4772_/B sky130_fd_sc_hd__a21o_1
X_6508_ _6466_/A _6493_/C _5721_/A _6507_/Y vssd1 vssd1 vccd1 vccd1 _6565_/A sky130_fd_sc_hd__o211a_1
X_6439_ _6439_/A _6439_/B vssd1 vssd1 vccd1 vccd1 _6441_/B sky130_fd_sc_hd__nor2_1
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold10 hold9/X vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_75_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold65/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__clkbuf_1
Xhold87 hold87/A vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_90_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_7 _5210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6790_ _6788_/X _6789_/Y _6261_/A vssd1 vssd1 vccd1 vccd1 _6790_/X sky130_fd_sc_hd__a21o_1
X_5810_ _5810_/A _6084_/A vssd1 vssd1 vccd1 vccd1 _5811_/B sky130_fd_sc_hd__xnor2_2
XFILLER_62_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5741_ _6625_/A _5756_/A vssd1 vssd1 vccd1 vccd1 _6054_/A sky130_fd_sc_hd__or2_2
X_7411_ _7411_/A _3707_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[15] sky130_fd_sc_hd__ebufn_8
X_5672_ _5722_/A _5873_/A _5694_/A vssd1 vssd1 vccd1 vccd1 _5673_/C sky130_fd_sc_hd__and3_1
XFILLER_30_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4623_ _4623_/A _4622_/B vssd1 vssd1 vccd1 vccd1 _4623_/X sky130_fd_sc_hd__or2b_1
X_4554_ _4554_/A _4554_/B vssd1 vssd1 vccd1 vccd1 _4652_/A sky130_fd_sc_hd__xnor2_1
X_7342_ _7342_/A _3626_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[16] sky130_fd_sc_hd__ebufn_8
XFILLER_89_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4485_ _4485_/A _4485_/B vssd1 vssd1 vccd1 vccd1 _4486_/B sky130_fd_sc_hd__or2_1
X_6224_ _6153_/A _6153_/B _6223_/X vssd1 vssd1 vccd1 vccd1 _6298_/B sky130_fd_sc_hd__a21o_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6155_ _6055_/A _6055_/B _6154_/Y vssd1 vssd1 vccd1 vccd1 _6236_/B sky130_fd_sc_hd__a21o_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6086_ _5810_/A _6084_/Y _6085_/X vssd1 vssd1 vccd1 vccd1 _6089_/A sky130_fd_sc_hd__a21oi_2
X_5106_ _5106_/A _5254_/B vssd1 vssd1 vccd1 vccd1 _5107_/B sky130_fd_sc_hd__xor2_2
X_5037_ _5037_/A _5037_/B vssd1 vssd1 vccd1 vccd1 _5183_/B sky130_fd_sc_hd__xnor2_1
XFILLER_38_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6988_ _7095_/A vssd1 vssd1 vccd1 vccd1 _7063_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5939_ _6061_/B _6409_/B vssd1 vssd1 vccd1 vccd1 _5953_/B sky130_fd_sc_hd__nand2_1
XFILLER_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4270_ _4466_/A _4377_/B _4124_/A vssd1 vssd1 vccd1 vccd1 _5707_/B sky130_fd_sc_hd__a21oi_4
XFILLER_97_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6911_ hold56/A _6893_/B _6894_/A hold25/A vssd1 vssd1 vccd1 vccd1 _6911_/X sky130_fd_sc_hd__a22o_1
XFILLER_47_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6842_ _6842_/A _6842_/B vssd1 vssd1 vccd1 vccd1 _6844_/A sky130_fd_sc_hd__and2_1
XFILLER_62_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3985_ _4694_/B vssd1 vssd1 vccd1 vccd1 _4638_/B sky130_fd_sc_hd__buf_2
XFILLER_22_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6773_ _6773_/A _6773_/B vssd1 vssd1 vccd1 vccd1 _6809_/A sky130_fd_sc_hd__xor2_2
X_5724_ _5725_/A _5724_/B vssd1 vssd1 vccd1 vccd1 _5762_/B sky130_fd_sc_hd__xnor2_1
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5655_ _6439_/A _6679_/B _6507_/B vssd1 vssd1 vccd1 vccd1 _6014_/B sky130_fd_sc_hd__a21oi_2
X_4606_ _4606_/A _4606_/B vssd1 vssd1 vccd1 vccd1 _4692_/A sky130_fd_sc_hd__xnor2_2
X_5586_ _5553_/A _5553_/B _5552_/A vssd1 vssd1 vccd1 vccd1 _5587_/B sky130_fd_sc_hd__a21oi_1
X_4537_ _4608_/A _4608_/B vssd1 vssd1 vccd1 vccd1 _4539_/B sky130_fd_sc_hd__and2b_1
XFILLER_89_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4468_ _4468_/A _4579_/A vssd1 vssd1 vccd1 vccd1 _4569_/A sky130_fd_sc_hd__nor2_1
XFILLER_89_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7187_ _7221_/CLK _7187_/D vssd1 vssd1 vccd1 vccd1 _7187_/Q sky130_fd_sc_hd__dfxtp_1
X_6207_ _6207_/A _6207_/B vssd1 vssd1 vccd1 vccd1 _6263_/B sky130_fd_sc_hd__xor2_4
X_4399_ _4392_/B _4531_/B _4180_/X vssd1 vssd1 vccd1 vccd1 _4401_/B sky130_fd_sc_hd__a21oi_1
X_6138_ _6142_/B vssd1 vssd1 vccd1 vccd1 _7003_/A sky130_fd_sc_hd__clkbuf_4
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6069_ _6070_/A _6070_/B _6070_/C vssd1 vssd1 vccd1 vccd1 _6167_/A sky130_fd_sc_hd__a21o_1
XFILLER_26_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7308__101 vssd1 vssd1 vccd1 vccd1 _7308__101/HI _7416_/A sky130_fd_sc_hd__conb_1
XFILLER_42_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3770_ _3770_/A _3770_/B vssd1 vssd1 vccd1 vccd1 _3770_/Y sky130_fd_sc_hd__nand2_1
X_5440_ _5547_/A _5547_/B vssd1 vssd1 vccd1 vccd1 _5442_/A sky130_fd_sc_hd__nor2_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5371_ _5371_/A _5371_/B vssd1 vssd1 vccd1 vccd1 _5380_/A sky130_fd_sc_hd__xnor2_1
X_7110_ hold94/X _7114_/B vssd1 vssd1 vccd1 vccd1 _7110_/X sky130_fd_sc_hd__or2_1
X_4322_ _3770_/A _4458_/B _4321_/X vssd1 vssd1 vccd1 vccd1 _4456_/A sky130_fd_sc_hd__a21bo_1
XFILLER_99_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4253_ _4253_/A _4254_/B vssd1 vssd1 vccd1 vccd1 _4500_/B sky130_fd_sc_hd__xnor2_1
X_7041_ _7041_/A _7059_/B vssd1 vssd1 vccd1 vccd1 _7041_/X sky130_fd_sc_hd__or2_1
X_4184_ _4182_/A _4182_/B _4183_/X vssd1 vssd1 vccd1 vccd1 _4243_/B sky130_fd_sc_hd__o21ai_4
XFILLER_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_7_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7221_/CLK
+ sky130_fd_sc_hd__clkbuf_2
X_6825_ _6983_/A _6825_/B vssd1 vssd1 vccd1 vccd1 _6856_/B sky130_fd_sc_hd__nor2_1
X_3968_ _7158_/Q vssd1 vssd1 vccd1 vccd1 _6445_/B sky130_fd_sc_hd__buf_2
X_6756_ _5113_/X hold128/X _6754_/X _6755_/Y _6405_/X vssd1 vssd1 vccd1 vccd1 hold42/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5707_ _5708_/B _5707_/B vssd1 vssd1 vccd1 vccd1 _5709_/A sky130_fd_sc_hd__and2b_1
X_3899_ _4533_/A vssd1 vssd1 vccd1 vccd1 _7041_/A sky130_fd_sc_hd__clkbuf_2
X_6687_ _6926_/A _6687_/B vssd1 vssd1 vccd1 vccd1 _6688_/B sky130_fd_sc_hd__and2b_1
XFILLER_12_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5638_ _5899_/A _6698_/A vssd1 vssd1 vccd1 vccd1 _5900_/A sky130_fd_sc_hd__nor2_1
XFILLER_88_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5569_ _5569_/A _5569_/B _5569_/C vssd1 vssd1 vccd1 vccd1 _5570_/B sky130_fd_sc_hd__and3_1
XFILLER_5_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4940_ _4940_/A _4940_/B vssd1 vssd1 vccd1 vccd1 _4940_/X sky130_fd_sc_hd__and2_1
X_4871_ _4822_/B _4822_/C _7038_/A vssd1 vssd1 vccd1 vccd1 _4872_/B sky130_fd_sc_hd__a21o_1
XFILLER_60_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3822_ _7199_/Q vssd1 vssd1 vccd1 vccd1 _4956_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6610_ _6643_/A _6643_/B _6609_/Y vssd1 vssd1 vccd1 vccd1 _6710_/A sky130_fd_sc_hd__o21a_1
XFILLER_32_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6541_ _6541_/A _6541_/B vssd1 vssd1 vccd1 vccd1 _6544_/A sky130_fd_sc_hd__nor2_1
X_3753_ _7189_/Q vssd1 vssd1 vccd1 vccd1 _6120_/B sky130_fd_sc_hd__clkbuf_4
X_3684_ _3684_/A vssd1 vssd1 vccd1 vccd1 _3684_/Y sky130_fd_sc_hd__inv_2
X_6472_ _6475_/D _6472_/B vssd1 vssd1 vccd1 vccd1 _6473_/B sky130_fd_sc_hd__nand2_1
X_5423_ _5423_/A _5423_/B vssd1 vssd1 vccd1 vccd1 _5444_/A sky130_fd_sc_hd__nor2_1
X_5354_ _5235_/B _5354_/B vssd1 vssd1 vccd1 vccd1 _5355_/B sky130_fd_sc_hd__and2b_1
X_4305_ _7176_/Q _5167_/A vssd1 vssd1 vccd1 vccd1 _4469_/B sky130_fd_sc_hd__nand2_1
X_5285_ _5285_/A _5285_/B vssd1 vssd1 vccd1 vccd1 _5295_/A sky130_fd_sc_hd__nor2_1
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4236_ _4236_/A _4236_/B vssd1 vssd1 vccd1 vccd1 _4491_/A sky130_fd_sc_hd__xor2_4
X_7024_ _6137_/B _7018_/X _7023_/X _7021_/X vssd1 vssd1 vccd1 vccd1 _7187_/D sky130_fd_sc_hd__o211a_1
XFILLER_101_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4167_ _4167_/A _4167_/B vssd1 vssd1 vccd1 vccd1 _5098_/A sky130_fd_sc_hd__xnor2_2
XFILLER_55_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4098_ _4225_/A vssd1 vssd1 vccd1 vccd1 _6761_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_70_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6808_ _6808_/A _6808_/B vssd1 vssd1 vccd1 vccd1 _6837_/A sky130_fd_sc_hd__xor2_1
XFILLER_23_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6739_ _6739_/A _6774_/A vssd1 vssd1 vccd1 vccd1 _6740_/B sky130_fd_sc_hd__xnor2_1
XFILLER_78_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5070_ _5218_/A _5220_/B vssd1 vssd1 vccd1 vccd1 _5071_/B sky130_fd_sc_hd__xor2_1
X_4021_ _3997_/B _4022_/A vssd1 vssd1 vccd1 vccd1 _4021_/X sky130_fd_sc_hd__and2b_1
XFILLER_1_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5972_ _6954_/A _6693_/A _5972_/C vssd1 vssd1 vccd1 vccd1 _5981_/A sky130_fd_sc_hd__nand3_1
XFILLER_52_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4923_ _4923_/A _4907_/A vssd1 vssd1 vccd1 vccd1 _4923_/X sky130_fd_sc_hd__or2b_1
XFILLER_18_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4854_ _4902_/A _4902_/B vssd1 vssd1 vccd1 vccd1 _4903_/A sky130_fd_sc_hd__nand2_1
XFILLER_33_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4785_ _4785_/A _4785_/B vssd1 vssd1 vccd1 vccd1 _4786_/A sky130_fd_sc_hd__nand2_1
X_3805_ _3805_/A _3805_/B vssd1 vssd1 vccd1 vccd1 _4481_/A sky130_fd_sc_hd__nand2_1
X_3736_ _3739_/A vssd1 vssd1 vccd1 vccd1 _3736_/Y sky130_fd_sc_hd__inv_2
X_6524_ _6524_/A _6524_/B vssd1 vssd1 vccd1 vccd1 _6524_/X sky130_fd_sc_hd__and2_1
X_6455_ _6455_/A _6455_/B vssd1 vssd1 vccd1 vccd1 _6458_/B sky130_fd_sc_hd__nand2_1
X_3667_ _3679_/A vssd1 vssd1 vccd1 vccd1 _3672_/A sky130_fd_sc_hd__buf_12
X_6386_ _6969_/A _6323_/B _6353_/B _6385_/X vssd1 vssd1 vccd1 vccd1 _6387_/B sky130_fd_sc_hd__a31oi_2
X_5406_ _5406_/A vssd1 vssd1 vccd1 vccd1 _6523_/A sky130_fd_sc_hd__buf_2
X_5337_ _5337_/A _5337_/B vssd1 vssd1 vccd1 vccd1 _5423_/B sky130_fd_sc_hd__xor2_2
X_5268_ _5275_/A vssd1 vssd1 vccd1 vccd1 _5391_/A sky130_fd_sc_hd__clkbuf_2
X_4219_ _4422_/A _4422_/B _4218_/Y vssd1 vssd1 vccd1 vccd1 _4220_/B sky130_fd_sc_hd__a21oi_1
XFILLER_75_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7007_ _7007_/A vssd1 vssd1 vccd1 vccd1 _7007_/X sky130_fd_sc_hd__buf_2
XFILLER_56_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5199_ _5199_/A _5199_/B vssd1 vssd1 vccd1 vccd1 _5430_/A sky130_fd_sc_hd__and2_1
XFILLER_55_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4570_ _4658_/A _4570_/B vssd1 vssd1 vccd1 vccd1 _4665_/B sky130_fd_sc_hd__xnor2_1
X_6240_ _6240_/A vssd1 vssd1 vccd1 vccd1 _6413_/A sky130_fd_sc_hd__clkbuf_2
X_6171_ _6171_/A _6171_/B vssd1 vssd1 vccd1 vccd1 _6171_/X sky130_fd_sc_hd__or2_1
XFILLER_97_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5122_ _7215_/Q _5122_/B _5277_/B vssd1 vssd1 vccd1 vccd1 _5124_/A sky130_fd_sc_hd__or3_1
X_5053_ _5190_/B _5053_/B vssd1 vssd1 vccd1 vccd1 _5054_/B sky130_fd_sc_hd__xnor2_2
XFILLER_84_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4004_ _4004_/A _4649_/A vssd1 vssd1 vccd1 vccd1 _4176_/B sky130_fd_sc_hd__and2_2
XFILLER_37_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5955_ _5955_/A _5955_/B vssd1 vssd1 vccd1 vccd1 _6001_/B sky130_fd_sc_hd__xnor2_1
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4906_ _4906_/A _4906_/B vssd1 vssd1 vccd1 vccd1 _4923_/A sky130_fd_sc_hd__nor2_1
X_5886_ _5886_/A _5886_/B vssd1 vssd1 vccd1 vccd1 _5887_/B sky130_fd_sc_hd__and2_1
X_4837_ _4837_/A _4837_/B vssd1 vssd1 vccd1 vccd1 _4838_/C sky130_fd_sc_hd__xor2_1
X_4768_ _7036_/A _4821_/B _4768_/C vssd1 vssd1 vccd1 vccd1 _4768_/X sky130_fd_sc_hd__and3_1
X_3719_ _3721_/A vssd1 vssd1 vccd1 vccd1 _3719_/Y sky130_fd_sc_hd__inv_2
X_4699_ _4763_/A _4697_/A _4763_/B _4698_/Y vssd1 vssd1 vccd1 vccd1 _4704_/B sky130_fd_sc_hd__o31a_1
X_6507_ _6507_/A _6507_/B vssd1 vssd1 vccd1 vccd1 _6507_/Y sky130_fd_sc_hd__nor2_1
X_6438_ _6470_/A _6455_/B vssd1 vssd1 vccd1 vccd1 _6443_/A sky130_fd_sc_hd__xnor2_2
X_6369_ _6852_/A _6369_/B vssd1 vssd1 vccd1 vccd1 _6370_/B sky130_fd_sc_hd__and2_1
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_48_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold77 hold77/A vssd1 vssd1 vccd1 vccd1 hold77/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold66 hold66/A vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_56_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_8 _5210_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5740_ _6136_/A _5718_/A _5714_/B _5714_/A vssd1 vssd1 vccd1 vccd1 _5744_/A sky130_fd_sc_hd__o22ai_2
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5671_ _6027_/A _5671_/B vssd1 vssd1 vccd1 vccd1 _5694_/A sky130_fd_sc_hd__xor2_4
X_7410_ _7410_/A _3706_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[14] sky130_fd_sc_hd__ebufn_8
X_4622_ _4623_/A _4622_/B vssd1 vssd1 vccd1 vccd1 _4690_/B sky130_fd_sc_hd__xnor2_1
XFILLER_30_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4553_ _4553_/A _4659_/B vssd1 vssd1 vccd1 vccd1 _4554_/B sky130_fd_sc_hd__nand2_1
X_7341_ _7341_/A _3622_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[15] sky130_fd_sc_hd__ebufn_8
X_7325__118 vssd1 vssd1 vccd1 vccd1 _7325__118/HI _7433_/A sky130_fd_sc_hd__conb_1
X_4484_ hold91/A _6624_/A _4785_/A vssd1 vssd1 vccd1 vccd1 _4485_/B sky130_fd_sc_hd__and3_1
X_6223_ _6150_/B _6223_/B vssd1 vssd1 vccd1 vccd1 _6223_/X sky130_fd_sc_hd__and2b_1
XFILLER_97_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6154_ _6154_/A _6154_/B vssd1 vssd1 vccd1 vccd1 _6154_/Y sky130_fd_sc_hd__nor2_1
XFILLER_97_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5105_ _4522_/A _4522_/B _5104_/X vssd1 vssd1 vccd1 vccd1 _5254_/B sky130_fd_sc_hd__a21bo_2
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6085_ _5800_/B _6085_/B vssd1 vssd1 vccd1 vccd1 _6085_/X sky130_fd_sc_hd__and2b_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5036_ _5036_/A _5036_/B vssd1 vssd1 vccd1 vccd1 _5037_/B sky130_fd_sc_hd__nor2_1
XFILLER_38_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6987_ _6828_/A _6977_/X _6986_/Y _6979_/X vssd1 vssd1 vccd1 vccd1 _7174_/D sky130_fd_sc_hd__o211a_1
X_5938_ _5938_/A _5938_/B vssd1 vssd1 vccd1 vccd1 _5953_/A sky130_fd_sc_hd__or2_1
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5869_ _5869_/A _5869_/B vssd1 vssd1 vccd1 vccd1 _5908_/A sky130_fd_sc_hd__xnor2_2
XFILLER_21_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7275__68 vssd1 vssd1 vccd1 vccd1 _7275__68/HI _7374_/A sky130_fd_sc_hd__conb_1
XFILLER_48_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6910_ _7116_/A hold12/X vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__nor2_1
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6841_ _6786_/A _6789_/Y _6840_/Y _6816_/B vssd1 vssd1 vccd1 vccd1 _6842_/B sky130_fd_sc_hd__a31o_1
X_3984_ _4526_/B _4873_/A vssd1 vssd1 vccd1 vccd1 _4694_/B sky130_fd_sc_hd__and2_1
XFILLER_22_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6772_ _6772_/A _6772_/B vssd1 vssd1 vccd1 vccd1 _6773_/B sky130_fd_sc_hd__xnor2_1
XFILLER_50_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5723_ _5723_/A _5723_/B vssd1 vssd1 vccd1 vccd1 _5724_/B sky130_fd_sc_hd__and2_2
X_5654_ _7153_/Q _5691_/B vssd1 vssd1 vccd1 vccd1 _6507_/B sky130_fd_sc_hd__nor2_2
XFILLER_30_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4605_ _4605_/A _4539_/X vssd1 vssd1 vccd1 vccd1 _4606_/A sky130_fd_sc_hd__or2b_1
XFILLER_30_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5585_ _5554_/A _5554_/B _5584_/Y vssd1 vssd1 vccd1 vccd1 _5587_/A sky130_fd_sc_hd__o21a_1
X_4536_ _7078_/A _4639_/B _4535_/Y vssd1 vssd1 vccd1 vccd1 _4608_/B sky130_fd_sc_hd__a21o_1
X_4467_ _5827_/A _4467_/B _4467_/C vssd1 vssd1 vccd1 vccd1 _4579_/A sky130_fd_sc_hd__and3_1
X_4398_ _7194_/Q _4531_/B vssd1 vssd1 vccd1 vccd1 _4401_/A sky130_fd_sc_hd__xnor2_1
X_7186_ _7221_/CLK _7186_/D vssd1 vssd1 vccd1 vccd1 _7186_/Q sky130_fd_sc_hd__dfxtp_2
X_6206_ _7053_/A _6206_/B vssd1 vssd1 vccd1 vccd1 _6207_/B sky130_fd_sc_hd__xnor2_2
X_6137_ _7006_/A _6137_/B vssd1 vssd1 vccd1 vccd1 _6145_/A sky130_fd_sc_hd__nor2_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6068_ _6228_/C _6068_/B vssd1 vssd1 vccd1 vccd1 _6070_/C sky130_fd_sc_hd__and2_1
XFILLER_38_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5019_ _5019_/A vssd1 vssd1 vccd1 vccd1 _5640_/A sky130_fd_sc_hd__buf_2
XFILLER_26_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5370_ _5468_/A _5468_/B vssd1 vssd1 vccd1 vccd1 _5371_/B sky130_fd_sc_hd__xnor2_2
X_4321_ _4321_/A _4320_/B vssd1 vssd1 vccd1 vccd1 _4321_/X sky130_fd_sc_hd__or2b_1
X_7040_ _7063_/A vssd1 vssd1 vccd1 vccd1 _7059_/B sky130_fd_sc_hd__clkbuf_1
X_4252_ _4252_/A _4506_/C vssd1 vssd1 vccd1 vccd1 _4254_/B sky130_fd_sc_hd__xnor2_1
X_4183_ _7083_/A _4394_/B vssd1 vssd1 vccd1 vccd1 _4183_/X sky130_fd_sc_hd__or2_1
XFILLER_79_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6824_ _6824_/A _6824_/B vssd1 vssd1 vccd1 vccd1 _6856_/A sky130_fd_sc_hd__nor2_1
XFILLER_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3967_ _3967_/A _3967_/B vssd1 vssd1 vccd1 vccd1 _5000_/B sky130_fd_sc_hd__nand2_1
X_6755_ _6751_/Y _6753_/Y _6752_/Y _5113_/X vssd1 vssd1 vccd1 vccd1 _6755_/Y sky130_fd_sc_hd__o31ai_1
X_5706_ _5715_/A _5706_/B vssd1 vssd1 vccd1 vccd1 _5708_/B sky130_fd_sc_hd__xnor2_1
X_3898_ _7194_/Q vssd1 vssd1 vccd1 vccd1 _4533_/A sky130_fd_sc_hd__clkbuf_2
X_6686_ _6698_/A _6698_/B _6684_/B _6685_/Y vssd1 vssd1 vccd1 vccd1 _6686_/X sky130_fd_sc_hd__a2bb2o_1
X_5637_ _5972_/C _5640_/A _6409_/A vssd1 vssd1 vccd1 vccd1 _6698_/A sky130_fd_sc_hd__mux2_2
X_5568_ _5569_/A _5569_/B _5569_/C vssd1 vssd1 vccd1 vccd1 _5570_/A sky130_fd_sc_hd__a21oi_1
X_4519_ _4520_/A _4520_/B vssd1 vssd1 vccd1 vccd1 _4599_/B sky130_fd_sc_hd__xor2_1
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5499_ _5499_/A _5499_/B vssd1 vssd1 vccd1 vccd1 _5513_/B sky130_fd_sc_hd__nor2_1
X_7169_ _7172_/CLK _7169_/D vssd1 vssd1 vccd1 vccd1 _7169_/Q sky130_fd_sc_hd__dfxtp_1
X_7245__38 vssd1 vssd1 vccd1 vccd1 _7245__38/HI _7344_/A sky130_fd_sc_hd__conb_1
XFILLER_85_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4870_ _4870_/A _4870_/B vssd1 vssd1 vccd1 vccd1 _4884_/A sky130_fd_sc_hd__xnor2_2
XFILLER_17_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3821_ _4426_/A vssd1 vssd1 vccd1 vccd1 _7089_/A sky130_fd_sc_hd__clkinv_2
XFILLER_20_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6540_ _6540_/A _6540_/B vssd1 vssd1 vccd1 vccd1 _6549_/A sky130_fd_sc_hd__or2_1
XFILLER_9_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3752_ _7099_/A vssd1 vssd1 vccd1 vccd1 _3752_/X sky130_fd_sc_hd__clkbuf_2
X_6471_ _6941_/A _6475_/B vssd1 vssd1 vccd1 vccd1 _6725_/A sky130_fd_sc_hd__nor2_1
X_3683_ _3684_/A vssd1 vssd1 vccd1 vccd1 _3683_/Y sky130_fd_sc_hd__inv_2
X_5422_ _5315_/A _5315_/B _5318_/B vssd1 vssd1 vccd1 vccd1 _5456_/A sky130_fd_sc_hd__a21bo_1
X_5353_ _5234_/A _5353_/B vssd1 vssd1 vccd1 vccd1 _5355_/A sky130_fd_sc_hd__and2b_1
X_4304_ _4304_/A _4304_/B vssd1 vssd1 vccd1 vccd1 _4338_/A sky130_fd_sc_hd__xnor2_2
XFILLER_99_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5284_ _5284_/A _5284_/B _5284_/C vssd1 vssd1 vccd1 vccd1 _5285_/B sky130_fd_sc_hd__nor3_1
XFILLER_101_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4235_ _4220_/A _4220_/B _4234_/X vssd1 vssd1 vccd1 vccd1 _4236_/B sky130_fd_sc_hd__o21a_4
X_7023_ _7023_/A _7025_/B vssd1 vssd1 vccd1 vccd1 _7023_/X sky130_fd_sc_hd__or2_1
X_4166_ _4166_/A _5045_/A vssd1 vssd1 vccd1 vccd1 _4167_/B sky130_fd_sc_hd__xnor2_1
X_4097_ _7166_/Q _4097_/B vssd1 vssd1 vccd1 vccd1 _4225_/A sky130_fd_sc_hd__xnor2_4
XFILLER_82_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6807_ _6833_/B _6807_/B vssd1 vssd1 vccd1 vccd1 _6808_/B sky130_fd_sc_hd__xnor2_1
X_4999_ _4150_/A _4150_/B _4164_/B _4163_/A vssd1 vssd1 vccd1 vccd1 _5037_/A sky130_fd_sc_hd__a31o_2
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6738_ _6536_/A _6536_/B _6737_/X vssd1 vssd1 vccd1 vccd1 _6774_/A sky130_fd_sc_hd__o21a_1
X_6669_ _6667_/A _6667_/B _6701_/A _6701_/B vssd1 vssd1 vccd1 vccd1 _6671_/B sky130_fd_sc_hd__o22a_1
XFILLER_48_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4020_ _4042_/B _4042_/A vssd1 vssd1 vccd1 vccd1 _4044_/A sky130_fd_sc_hd__and2b_1
X_5971_ _6954_/A _6693_/A _5972_/C vssd1 vssd1 vccd1 vccd1 _5971_/X sky130_fd_sc_hd__and3_1
XFILLER_25_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4922_ _4903_/A _4907_/X _4921_/Y _4906_/B vssd1 vssd1 vccd1 vccd1 _4922_/X sky130_fd_sc_hd__a211o_1
XFILLER_33_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4853_ _5812_/A _4746_/B _4852_/Y vssd1 vssd1 vccd1 vccd1 _4902_/B sky130_fd_sc_hd__a21bo_1
X_4784_ _4784_/A _4784_/B vssd1 vssd1 vccd1 vccd1 _4787_/A sky130_fd_sc_hd__xor2_1
X_3804_ _5737_/A _4789_/B vssd1 vssd1 vccd1 vccd1 _3805_/B sky130_fd_sc_hd__or2_1
X_3735_ _3739_/A vssd1 vssd1 vccd1 vccd1 _3735_/Y sky130_fd_sc_hd__inv_2
X_6523_ _6523_/A _6524_/B vssd1 vssd1 vccd1 vccd1 _6531_/B sky130_fd_sc_hd__xor2_1
X_6454_ _6454_/A _6454_/B vssd1 vssd1 vccd1 vccd1 _6458_/A sky130_fd_sc_hd__or2_1
XFILLER_9_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3666_ _3666_/A vssd1 vssd1 vccd1 vccd1 _3666_/Y sky130_fd_sc_hd__inv_2
X_5405_ _7096_/A _5293_/B _5294_/A _5290_/A vssd1 vssd1 vccd1 vccd1 _5500_/B sky130_fd_sc_hd__a31o_1
X_6385_ _6352_/B _6385_/B vssd1 vssd1 vccd1 vccd1 _6385_/X sky130_fd_sc_hd__and2b_1
XFILLER_87_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5336_ hold84/A _5335_/A _5210_/B _5335_/Y vssd1 vssd1 vccd1 vccd1 _5337_/B sky130_fd_sc_hd__a31o_1
X_5267_ _5267_/A _5267_/B vssd1 vssd1 vccd1 vccd1 _5271_/A sky130_fd_sc_hd__nand2_1
X_4218_ _4218_/A _4218_/B vssd1 vssd1 vccd1 vccd1 _4218_/Y sky130_fd_sc_hd__nor2_1
XFILLER_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7006_ _7006_/A _7006_/B vssd1 vssd1 vccd1 vccd1 _7006_/Y sky130_fd_sc_hd__nand2_1
XFILLER_18_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5198_ _7173_/Q _5198_/B vssd1 vssd1 vccd1 vccd1 _5199_/B sky130_fd_sc_hd__or2_1
XFILLER_68_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4149_ _4149_/A _4149_/B vssd1 vssd1 vccd1 vccd1 _4150_/B sky130_fd_sc_hd__or2_1
XFILLER_28_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6170_ _6170_/A _6170_/B vssd1 vssd1 vccd1 vccd1 _6173_/A sky130_fd_sc_hd__xor2_4
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5121_ _5121_/A vssd1 vssd1 vccd1 vccd1 _5122_/B sky130_fd_sc_hd__inv_2
XFILLER_97_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5052_ _3783_/A _5048_/A _5190_/A vssd1 vssd1 vccd1 vccd1 _5053_/B sky130_fd_sc_hd__a21oi_1
XFILLER_38_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4003_ _4003_/A _7208_/Q vssd1 vssd1 vccd1 vccd1 _4649_/A sky130_fd_sc_hd__or2b_1
XFILLER_77_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5954_ _5954_/A _5954_/B vssd1 vssd1 vccd1 vccd1 _6001_/A sky130_fd_sc_hd__nor2_1
X_4905_ _4905_/A _4905_/B vssd1 vssd1 vccd1 vccd1 _4906_/B sky130_fd_sc_hd__and2_1
X_5885_ _5886_/A _5886_/B vssd1 vssd1 vccd1 vccd1 _5887_/A sky130_fd_sc_hd__nor2_1
XFILLER_33_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4836_ _4836_/A vssd1 vssd1 vccd1 vccd1 _4836_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4767_ _4821_/A vssd1 vssd1 vccd1 vccd1 _7036_/A sky130_fd_sc_hd__clkbuf_2
X_6506_ _6506_/A _6506_/B _6506_/C vssd1 vssd1 vccd1 vccd1 _6541_/A sky130_fd_sc_hd__and3_1
X_4698_ _4761_/A _4761_/B vssd1 vssd1 vccd1 vccd1 _4698_/Y sky130_fd_sc_hd__nand2_1
X_3718_ _3721_/A vssd1 vssd1 vccd1 vccd1 _3718_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3649_ _3653_/A vssd1 vssd1 vccd1 vccd1 _3649_/Y sky130_fd_sc_hd__inv_2
X_6437_ _6454_/A _6441_/A vssd1 vssd1 vccd1 vccd1 _6455_/B sky130_fd_sc_hd__xnor2_2
X_6368_ _6528_/A vssd1 vssd1 vccd1 vccd1 _6852_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5319_ _5383_/A _5383_/B vssd1 vssd1 vccd1 vccd1 _5321_/C sky130_fd_sc_hd__xor2_1
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_6299_ _6235_/A _6235_/B _6298_/Y vssd1 vssd1 vccd1 vccd1 _6349_/B sky130_fd_sc_hd__a21bo_1
XFILLER_48_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold56/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold67 hold67/A vssd1 vssd1 vccd1 vccd1 hold67/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_45_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_9 _6966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5670_ _5669_/A _5669_/B _5669_/C vssd1 vssd1 vccd1 vccd1 _5673_/B sky130_fd_sc_hd__o21ai_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4621_ _4692_/A _4692_/B _4620_/X vssd1 vssd1 vccd1 vccd1 _4622_/B sky130_fd_sc_hd__a21bo_1
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7340_ _7340_/A _3621_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[14] sky130_fd_sc_hd__ebufn_8
X_4552_ hold80/A _4659_/A _4552_/C vssd1 vssd1 vccd1 vccd1 _4659_/B sky130_fd_sc_hd__nor3_1
X_4483_ _4595_/A vssd1 vssd1 vccd1 vccd1 _4785_/A sky130_fd_sc_hd__inv_2
X_6222_ _6283_/A _6222_/B vssd1 vssd1 vccd1 vccd1 _6298_/A sky130_fd_sc_hd__xnor2_4
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6153_ _6153_/A _6153_/B vssd1 vssd1 vccd1 vccd1 _6156_/A sky130_fd_sc_hd__xnor2_4
XFILLER_97_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5104_ _5104_/A _4525_/A vssd1 vssd1 vccd1 vccd1 _5104_/X sky130_fd_sc_hd__or2b_1
XFILLER_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6084_ _6084_/A vssd1 vssd1 vccd1 vccd1 _6084_/Y sky130_fd_sc_hd__inv_2
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5035_ _5035_/A _5035_/B _5035_/C vssd1 vssd1 vccd1 vccd1 _5036_/B sky130_fd_sc_hd__nor3_1
X_6986_ _6986_/A _7006_/B vssd1 vssd1 vccd1 vccd1 _6986_/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5937_ _6160_/A _5937_/B vssd1 vssd1 vccd1 vccd1 _5938_/B sky130_fd_sc_hd__and2b_1
XFILLER_25_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5868_ _5868_/A _5868_/B vssd1 vssd1 vccd1 vccd1 _5886_/A sky130_fd_sc_hd__xnor2_1
X_4819_ _4819_/A _4819_/B vssd1 vssd1 vccd1 vccd1 _4870_/A sky130_fd_sc_hd__and2_1
XFILLER_31_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5799_ _6076_/B _5799_/B vssd1 vssd1 vccd1 vccd1 _5800_/B sky130_fd_sc_hd__or2_1
XFILLER_5_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6840_ _6840_/A vssd1 vssd1 vccd1 vccd1 _6840_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6771_ _6981_/A _6771_/B vssd1 vssd1 vccd1 vccd1 _6772_/B sky130_fd_sc_hd__xnor2_1
X_5722_ _5722_/A _5873_/A vssd1 vssd1 vccd1 vccd1 _5723_/B sky130_fd_sc_hd__or2_1
X_3983_ _3983_/A _3983_/B vssd1 vssd1 vccd1 vccd1 _4045_/A sky130_fd_sc_hd__xor2_1
XFILLER_62_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5653_ _6434_/A vssd1 vssd1 vccd1 vccd1 _6679_/B sky130_fd_sc_hd__buf_2
X_4604_ _4604_/A _4604_/B vssd1 vssd1 vccd1 vccd1 _4623_/A sky130_fd_sc_hd__xnor2_2
X_5584_ _5584_/A _5584_/B vssd1 vssd1 vccd1 vccd1 _5584_/Y sky130_fd_sc_hd__nand2_1
X_4535_ _4535_/A _4766_/A vssd1 vssd1 vccd1 vccd1 _4535_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4466_ _4466_/A _4745_/B vssd1 vssd1 vccd1 vccd1 _4467_/C sky130_fd_sc_hd__or2_1
X_4397_ _4505_/A _4397_/B vssd1 vssd1 vccd1 vccd1 _4498_/A sky130_fd_sc_hd__xor2_2
X_7185_ _7225_/CLK _7185_/D vssd1 vssd1 vccd1 vccd1 _7185_/Q sky130_fd_sc_hd__dfxtp_4
X_6205_ _6118_/A _6118_/B _6122_/B _6125_/A vssd1 vssd1 vccd1 vccd1 _6207_/A sky130_fd_sc_hd__a31o_1
XFILLER_58_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6136_ _6136_/A vssd1 vssd1 vccd1 vccd1 _7006_/A sky130_fd_sc_hd__clkbuf_2
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6067_ _6067_/A _6286_/B vssd1 vssd1 vccd1 vccd1 _6068_/B sky130_fd_sc_hd__or2_1
XFILLER_85_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5018_ _7114_/A _6941_/A _4154_/B _5017_/X vssd1 vssd1 vccd1 vccd1 _5174_/B sky130_fd_sc_hd__a31o_1
XFILLER_38_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6969_ _6969_/A _6975_/B vssd1 vssd1 vccd1 vccd1 _6969_/X sky130_fd_sc_hd__or2_1
XFILLER_13_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4320_ _4321_/A _4320_/B vssd1 vssd1 vccd1 vccd1 _4458_/B sky130_fd_sc_hd__xnor2_1
X_4251_ _4502_/A _4763_/A _4009_/B vssd1 vssd1 vccd1 vccd1 _4253_/A sky130_fd_sc_hd__o21a_1
XFILLER_95_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4182_ _4182_/A _4182_/B vssd1 vssd1 vccd1 vccd1 _4394_/B sky130_fd_sc_hd__xnor2_1
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6823_ _6986_/A _6852_/B vssd1 vssd1 vccd1 vccd1 _6827_/A sky130_fd_sc_hd__xnor2_1
XFILLER_35_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3966_ _3966_/A _3918_/A vssd1 vssd1 vccd1 vccd1 _3967_/B sky130_fd_sc_hd__or2b_1
XFILLER_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6754_ _6751_/Y _6752_/Y _6753_/Y vssd1 vssd1 vccd1 vccd1 _6754_/X sky130_fd_sc_hd__o21a_1
X_6685_ _6685_/A vssd1 vssd1 vccd1 vccd1 _6685_/Y sky130_fd_sc_hd__clkinv_2
X_5705_ _6142_/B hold89/A vssd1 vssd1 vccd1 vccd1 _5706_/B sky130_fd_sc_hd__xnor2_1
X_3897_ _3904_/A _3905_/B vssd1 vssd1 vccd1 vccd1 _3921_/A sky130_fd_sc_hd__xnor2_1
X_5636_ _5636_/A _5636_/B vssd1 vssd1 vccd1 vccd1 _5899_/A sky130_fd_sc_hd__or2_1
X_5567_ _5567_/A _5567_/B vssd1 vssd1 vccd1 vccd1 _5569_/C sky130_fd_sc_hd__xor2_1
X_4518_ _4601_/A _4601_/B _4517_/X vssd1 vssd1 vccd1 vccd1 _4520_/B sky130_fd_sc_hd__a21oi_1
Xhold120 _7036_/A vssd1 vssd1 vccd1 vccd1 hold120/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_5498_ _5498_/A _5498_/B vssd1 vssd1 vccd1 vccd1 _5513_/A sky130_fd_sc_hd__and2_1
X_4449_ _4795_/B vssd1 vssd1 vccd1 vccd1 _5644_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_77_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7168_ _7172_/CLK _7168_/D vssd1 vssd1 vccd1 vccd1 _7168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7099_ _7099_/A vssd1 vssd1 vccd1 vccd1 _7099_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6119_ _6120_/A _7025_/A _6120_/B vssd1 vssd1 vccd1 vccd1 _6121_/A sky130_fd_sc_hd__a21oi_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3820_ _7212_/Q vssd1 vssd1 vccd1 vccd1 _4426_/A sky130_fd_sc_hd__buf_2
XFILLER_60_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3751_ _7020_/A vssd1 vssd1 vccd1 vccd1 _7099_/A sky130_fd_sc_hd__buf_2
XFILLER_32_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6470_ _6470_/A _6943_/A vssd1 vssd1 vccd1 vccd1 _6475_/B sky130_fd_sc_hd__nand2_1
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3682_ _3684_/A vssd1 vssd1 vccd1 vccd1 _3682_/Y sky130_fd_sc_hd__inv_2
X_5421_ _5356_/A _5356_/B _5420_/X vssd1 vssd1 vccd1 vccd1 _5457_/A sky130_fd_sc_hd__o21ai_1
X_5352_ _5352_/A _5352_/B vssd1 vssd1 vccd1 vccd1 _5356_/A sky130_fd_sc_hd__xnor2_2
X_4303_ _4303_/A _4385_/B vssd1 vssd1 vccd1 vccd1 _4304_/B sky130_fd_sc_hd__xnor2_2
XFILLER_101_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7022_ hold89/X _7018_/X _7019_/X _7021_/X vssd1 vssd1 vccd1 vccd1 _7186_/D sky130_fd_sc_hd__o211a_1
X_5283_ _5284_/A _5284_/B _5284_/C vssd1 vssd1 vccd1 vccd1 _5285_/A sky130_fd_sc_hd__o21a_1
XFILLER_101_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4234_ _4421_/A _4421_/B vssd1 vssd1 vccd1 vccd1 _4234_/X sky130_fd_sc_hd__or2b_1
XFILLER_4_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4165_ _4165_/A _4165_/B vssd1 vssd1 vccd1 vccd1 _5045_/A sky130_fd_sc_hd__xnor2_1
XFILLER_95_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4096_ _5002_/A _4096_/B vssd1 vssd1 vccd1 vccd1 _4372_/A sky130_fd_sc_hd__xnor2_2
XFILLER_51_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6806_ _6772_/A _6772_/B _6773_/B _6773_/A vssd1 vssd1 vccd1 vccd1 _6807_/B sky130_fd_sc_hd__o2bb2a_1
X_4998_ _4998_/A _4998_/B vssd1 vssd1 vccd1 vccd1 _5183_/A sky130_fd_sc_hd__xnor2_1
XFILLER_11_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3949_ _3963_/A _3963_/B vssd1 vssd1 vccd1 vccd1 _4024_/A sky130_fd_sc_hd__xnor2_2
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6737_ _6737_/A _6535_/B vssd1 vssd1 vccd1 vccd1 _6737_/X sky130_fd_sc_hd__or2b_1
X_6668_ _6241_/A _5796_/B _6668_/S vssd1 vssd1 vccd1 vccd1 _6701_/B sky130_fd_sc_hd__mux2_1
X_6599_ _6597_/A _6597_/B _6635_/A vssd1 vssd1 vccd1 vccd1 _6603_/B sky130_fd_sc_hd__o21ba_1
X_5619_ _5625_/A _5619_/B vssd1 vssd1 vccd1 vccd1 _5737_/C sky130_fd_sc_hd__or2_1
X_7305__98 vssd1 vssd1 vccd1 vccd1 _7305__98/HI _7413_/A sky130_fd_sc_hd__conb_1
XFILLER_2_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5970_ _6409_/A vssd1 vssd1 vccd1 vccd1 _6954_/A sky130_fd_sc_hd__buf_2
XFILLER_92_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4921_ _4905_/A _4905_/B _4913_/X _5911_/A _4920_/X vssd1 vssd1 vccd1 vccd1 _4921_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_64_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4852_ _6999_/A _5880_/B vssd1 vssd1 vccd1 vccd1 _4852_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3803_ _7171_/Q vssd1 vssd1 vccd1 vccd1 _5737_/A sky130_fd_sc_hd__clkbuf_2
X_4783_ _4788_/A _4788_/B _4782_/Y vssd1 vssd1 vccd1 vccd1 _4784_/B sky130_fd_sc_hd__a21oi_1
X_6522_ _6522_/A _6522_/B vssd1 vssd1 vccd1 vccd1 _6524_/B sky130_fd_sc_hd__xnor2_2
X_3734_ _3734_/A vssd1 vssd1 vccd1 vccd1 _3739_/A sky130_fd_sc_hd__buf_12
X_6453_ _6453_/A _6453_/B vssd1 vssd1 vccd1 vccd1 _6727_/A sky130_fd_sc_hd__or2_1
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3665_ _3666_/A vssd1 vssd1 vccd1 vccd1 _3665_/Y sky130_fd_sc_hd__inv_2
X_5404_ _5308_/B _5314_/B _5308_/A vssd1 vssd1 vccd1 vccd1 _5415_/A sky130_fd_sc_hd__o21ba_1
X_6384_ _6874_/A vssd1 vssd1 vccd1 vccd1 _6969_/A sky130_fd_sc_hd__buf_2
X_5335_ _5335_/A _5335_/B vssd1 vssd1 vccd1 vccd1 _5335_/Y sky130_fd_sc_hd__nor2_1
X_5266_ _5266_/A _5266_/B _5289_/B vssd1 vssd1 vccd1 vccd1 _5284_/B sky130_fd_sc_hd__and3_1
X_7005_ _7045_/A vssd1 vssd1 vccd1 vccd1 _7005_/X sky130_fd_sc_hd__buf_2
X_4217_ _4218_/A _4218_/B vssd1 vssd1 vccd1 vccd1 _4422_/B sky130_fd_sc_hd__xor2_2
XFILLER_68_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5197_ _6802_/A _6537_/B vssd1 vssd1 vccd1 vccd1 _5333_/A sky130_fd_sc_hd__or2_2
X_4148_ _4149_/A _4149_/B vssd1 vssd1 vccd1 vccd1 _4150_/A sky130_fd_sc_hd__nand2_1
X_4079_ _4197_/A _4080_/B vssd1 vssd1 vccd1 vccd1 _4204_/B sky130_fd_sc_hd__xnor2_1
XFILLER_70_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5120_ _5120_/A _5120_/B vssd1 vssd1 vccd1 vccd1 _5127_/B sky130_fd_sc_hd__nor2_1
XFILLER_69_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7296__89 vssd1 vssd1 vccd1 vccd1 _7296__89/HI _7404_/A sky130_fd_sc_hd__conb_1
X_5051_ _5051_/A vssd1 vssd1 vccd1 vccd1 _5190_/B sky130_fd_sc_hd__inv_2
X_4002_ _4002_/A _4002_/B vssd1 vssd1 vccd1 vccd1 _4176_/A sky130_fd_sc_hd__xnor2_1
XFILLER_65_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5953_ _5953_/A _5953_/B vssd1 vssd1 vccd1 vccd1 _5954_/B sky130_fd_sc_hd__and2_1
XFILLER_52_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4904_ _4904_/A _4904_/B vssd1 vssd1 vccd1 vccd1 _4905_/B sky130_fd_sc_hd__xnor2_1
X_5884_ _5908_/A _5908_/B _5883_/Y vssd1 vssd1 vccd1 vccd1 _5886_/B sky130_fd_sc_hd__a21oi_1
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4835_ _4837_/A _4837_/B vssd1 vssd1 vccd1 vccd1 _4836_/A sky130_fd_sc_hd__nor2_1
X_4766_ _4766_/A _4766_/B vssd1 vssd1 vccd1 vccd1 _4820_/B sky130_fd_sc_hd__and2_1
X_3717_ _3721_/A vssd1 vssd1 vccd1 vccd1 _3717_/Y sky130_fd_sc_hd__inv_2
X_6505_ _6505_/A _6505_/B _6505_/C vssd1 vssd1 vccd1 vccd1 _6506_/C sky130_fd_sc_hd__and3_1
X_4697_ _4697_/A _4697_/B vssd1 vssd1 vccd1 vccd1 _4761_/B sky130_fd_sc_hd__xnor2_2
X_3648_ _3648_/A vssd1 vssd1 vccd1 vccd1 _3653_/A sky130_fd_sc_hd__buf_12
X_6436_ _6454_/B vssd1 vssd1 vccd1 vccd1 _6441_/A sky130_fd_sc_hd__inv_2
X_6367_ _6824_/A vssd1 vssd1 vccd1 vccd1 _6990_/A sky130_fd_sc_hd__buf_2
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5318_ _5318_/A _5318_/B vssd1 vssd1 vccd1 vccd1 _5383_/B sky130_fd_sc_hd__nand2_1
X_6298_ _6298_/A _6298_/B vssd1 vssd1 vccd1 vccd1 _6298_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5249_ _5249_/A _5249_/B vssd1 vssd1 vccd1 vccd1 _5372_/A sky130_fd_sc_hd__xor2_4
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold68 hold68/A vssd1 vssd1 vccd1 vccd1 hold68/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_28_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4620_ _4620_/A _4619_/A vssd1 vssd1 vccd1 vccd1 _4620_/X sky130_fd_sc_hd__or2b_1
X_4551_ hold77/A _6439_/B vssd1 vssd1 vccd1 vccd1 _4552_/C sky130_fd_sc_hd__and2b_1
X_4482_ _4485_/A _4482_/B vssd1 vssd1 vccd1 vccd1 _4595_/A sky130_fd_sc_hd__or2_2
X_6221_ _6983_/A _6290_/B vssd1 vssd1 vccd1 vccd1 _6222_/B sky130_fd_sc_hd__xnor2_2
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6152_ _6575_/A _6226_/B vssd1 vssd1 vccd1 vccd1 _6153_/B sky130_fd_sc_hd__xor2_4
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ _5250_/A _5250_/B vssd1 vssd1 vccd1 vccd1 _5106_/A sky130_fd_sc_hd__xnor2_4
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ _6954_/A _5850_/B _5857_/B _5856_/A vssd1 vssd1 vccd1 vccd1 _6090_/A sky130_fd_sc_hd__a31o_2
XFILLER_85_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _5035_/A _5035_/B _5035_/C vssd1 vssd1 vccd1 vccd1 _5036_/A sky130_fd_sc_hd__o21a_1
XFILLER_53_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6985_ _7080_/A vssd1 vssd1 vccd1 vccd1 _7006_/B sky130_fd_sc_hd__clkbuf_4
X_5936_ _5936_/A vssd1 vssd1 vccd1 vccd1 _6947_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5867_ _5867_/A _5867_/B vssd1 vssd1 vccd1 vccd1 _5907_/A sky130_fd_sc_hd__and2_1
X_4818_ _4802_/A _4802_/C _4802_/B vssd1 vssd1 vccd1 vccd1 _4819_/B sky130_fd_sc_hd__o21ai_1
X_5798_ _5798_/A _5798_/B vssd1 vssd1 vccd1 vccd1 _5799_/B sky130_fd_sc_hd__and2_1
X_4749_ _4789_/B vssd1 vssd1 vccd1 vccd1 _6687_/B sky130_fd_sc_hd__clkbuf_2
X_6419_ _6627_/A vssd1 vssd1 vccd1 vccd1 _6679_/A sky130_fd_sc_hd__buf_2
X_7399_ _7399_/A _3693_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[3] sky130_fd_sc_hd__ebufn_8
XFILLER_48_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7266__59 vssd1 vssd1 vccd1 vccd1 _7266__59/HI _7365_/A sky130_fd_sc_hd__conb_1
XFILLER_94_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3982_ _3982_/A _5001_/B vssd1 vssd1 vccd1 vccd1 _3983_/B sky130_fd_sc_hd__xnor2_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6770_ _6802_/A _6802_/B vssd1 vssd1 vccd1 vccd1 _6771_/B sky130_fd_sc_hd__xnor2_1
X_5721_ _5721_/A _5721_/B vssd1 vssd1 vccd1 vccd1 _5725_/A sky130_fd_sc_hd__nand2_1
XFILLER_50_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5652_ _7153_/Q _7152_/Q vssd1 vssd1 vccd1 vccd1 _6434_/A sky130_fd_sc_hd__xor2_1
X_4603_ _4603_/A _4603_/B vssd1 vssd1 vccd1 vccd1 _4690_/A sky130_fd_sc_hd__nor2_1
X_5583_ _5557_/A _5578_/X _5581_/Y _5582_/Y vssd1 vssd1 vccd1 vccd1 _5588_/A sky130_fd_sc_hd__o31a_1
X_4534_ _4535_/A _4766_/A vssd1 vssd1 vccd1 vccd1 _4639_/B sky130_fd_sc_hd__xor2_1
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4465_ _4466_/A _4465_/B vssd1 vssd1 vccd1 vccd1 _4467_/B sky130_fd_sc_hd__nand2_1
X_4396_ _4504_/A _4504_/B vssd1 vssd1 vccd1 vccd1 _4505_/A sky130_fd_sc_hd__nor2_1
XFILLER_89_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7184_ _7225_/CLK _7184_/D vssd1 vssd1 vccd1 vccd1 _7184_/Q sky130_fd_sc_hd__dfxtp_2
X_6204_ _6204_/A _6204_/B vssd1 vssd1 vccd1 vccd1 _6263_/A sky130_fd_sc_hd__xnor2_4
XFILLER_97_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6135_ _6217_/A _6217_/B vssd1 vssd1 vccd1 vccd1 _6146_/A sky130_fd_sc_hd__xnor2_2
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6066_ _6067_/A _6286_/B vssd1 vssd1 vccd1 vccd1 _6228_/C sky130_fd_sc_hd__nand2_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5017_ _5017_/A _5017_/B vssd1 vssd1 vccd1 vccd1 _5017_/X sky130_fd_sc_hd__and2_1
XFILLER_45_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7280__73 vssd1 vssd1 vccd1 vccd1 _7280__73/HI _7379_/A sky130_fd_sc_hd__conb_1
X_6968_ _6943_/A _6964_/X _6966_/Y _6967_/X vssd1 vssd1 vccd1 vccd1 _7166_/D sky130_fd_sc_hd__o211a_1
X_5919_ _5950_/A _5950_/B vssd1 vssd1 vccd1 vccd1 _5919_/X sky130_fd_sc_hd__or2b_1
X_6899_ hold32/X _6890_/X _6898_/X vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__a21oi_1
XFILLER_42_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7315__108 vssd1 vssd1 vccd1 vccd1 _7315__108/HI _7423_/A sky130_fd_sc_hd__conb_1
XFILLER_76_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4250_ _4613_/A _5671_/B vssd1 vssd1 vccd1 vccd1 _4763_/A sky130_fd_sc_hd__xnor2_4
XFILLER_101_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4181_ _4533_/A _4531_/B _4180_/X vssd1 vssd1 vccd1 vccd1 _4182_/B sky130_fd_sc_hd__a21oi_2
XFILLER_86_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6822_ _6824_/A _6851_/B vssd1 vssd1 vccd1 vccd1 _6852_/B sky130_fd_sc_hd__xnor2_1
XFILLER_90_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3965_ _3965_/A _3909_/B vssd1 vssd1 vccd1 vccd1 _3967_/A sky130_fd_sc_hd__or2b_1
X_6753_ _6647_/A _6647_/B _6707_/A _6707_/B vssd1 vssd1 vccd1 vccd1 _6753_/Y sky130_fd_sc_hd__o22ai_4
X_3896_ _3896_/A _3896_/B vssd1 vssd1 vccd1 vccd1 _3905_/B sky130_fd_sc_hd__nand2_1
X_6684_ _6685_/A _6684_/B vssd1 vssd1 vccd1 vccd1 _6698_/B sky130_fd_sc_hd__xor2_1
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5704_ _5717_/A vssd1 vssd1 vccd1 vccd1 _6142_/B sky130_fd_sc_hd__clkbuf_2
X_5635_ _6571_/A _6589_/A _5611_/C vssd1 vssd1 vccd1 vccd1 _5636_/B sky130_fd_sc_hd__a21oi_1
Xhold110 _7109_/X vssd1 vssd1 vccd1 vccd1 _7220_/D sky130_fd_sc_hd__clkdlybuf4s50_1
X_5566_ _5526_/A _5526_/B _5525_/A vssd1 vssd1 vccd1 vccd1 _5567_/B sky130_fd_sc_hd__a21o_1
X_4517_ _4516_/A _4517_/B vssd1 vssd1 vccd1 vccd1 _4517_/X sky130_fd_sc_hd__and2b_1
Xhold121 _7023_/A vssd1 vssd1 vccd1 vccd1 hold121/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5497_ _5556_/A _5497_/B vssd1 vssd1 vccd1 vccd1 _5515_/A sky130_fd_sc_hd__or2_1
X_4448_ _7160_/Q vssd1 vssd1 vccd1 vccd1 _4795_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7167_ _7183_/CLK _7167_/D vssd1 vssd1 vccd1 vccd1 _7167_/Q sky130_fd_sc_hd__dfxtp_1
X_4379_ _4379_/A _4379_/B vssd1 vssd1 vccd1 vccd1 _5076_/A sky130_fd_sc_hd__xnor2_1
X_7098_ hold80/X _7106_/B vssd1 vssd1 vccd1 vccd1 hold81/A sky130_fd_sc_hd__or2_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6118_ _6118_/A _6118_/B vssd1 vssd1 vccd1 vccd1 _6122_/A sky130_fd_sc_hd__nand2_1
XFILLER_58_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6049_ _6049_/A _6049_/B vssd1 vssd1 vccd1 vccd1 _6049_/Y sky130_fd_sc_hd__nor2_1
XFILLER_37_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7236__29 vssd1 vssd1 vccd1 vccd1 _7236__29/HI _7335_/A sky130_fd_sc_hd__conb_1
XFILLER_76_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3750_ _5594_/A vssd1 vssd1 vccd1 vccd1 _3750_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3681_ _3684_/A vssd1 vssd1 vccd1 vccd1 _3681_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5420_ _5420_/A _5357_/B vssd1 vssd1 vccd1 vccd1 _5420_/X sky130_fd_sc_hd__or2b_1
X_5351_ _5351_/A _5351_/B vssd1 vssd1 vccd1 vccd1 _5352_/B sky130_fd_sc_hd__and2_1
XFILLER_99_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5282_ _5282_/A _5384_/B vssd1 vssd1 vccd1 vccd1 _5284_/C sky130_fd_sc_hd__xnor2_1
X_4302_ _4370_/A _4370_/B vssd1 vssd1 vccd1 vccd1 _4385_/B sky130_fd_sc_hd__xor2_2
X_7021_ _7073_/A vssd1 vssd1 vccd1 vccd1 _7021_/X sky130_fd_sc_hd__clkbuf_2
X_4233_ _4293_/A _4233_/B vssd1 vssd1 vccd1 vccd1 _4421_/B sky130_fd_sc_hd__xnor2_4
XFILLER_67_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4164_ _4164_/A _4164_/B vssd1 vssd1 vccd1 vccd1 _4165_/B sky130_fd_sc_hd__xnor2_4
XFILLER_83_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4095_ _4573_/A _4092_/Y _4094_/Y vssd1 vssd1 vccd1 vccd1 _4096_/B sky130_fd_sc_hd__o21a_1
XFILLER_55_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7250__43 vssd1 vssd1 vccd1 vccd1 _7250__43/HI _7349_/A sky130_fd_sc_hd__conb_1
XFILLER_36_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6805_ _6805_/A _6805_/B vssd1 vssd1 vccd1 vccd1 _6833_/B sky130_fd_sc_hd__xor2_1
X_4997_ _3983_/A _3983_/B _4996_/X vssd1 vssd1 vccd1 vccd1 _4998_/B sky130_fd_sc_hd__a21oi_2
XFILLER_11_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6736_ _6736_/A _6736_/B vssd1 vssd1 vccd1 vccd1 _6739_/A sky130_fd_sc_hd__xnor2_2
X_3948_ _4026_/A _4026_/B _3947_/Y vssd1 vssd1 vccd1 vccd1 _3963_/B sky130_fd_sc_hd__a21oi_1
X_6667_ _6667_/A _6667_/B vssd1 vssd1 vccd1 vccd1 _6701_/A sky130_fd_sc_hd__xnor2_1
X_3879_ _7093_/A _3879_/B vssd1 vssd1 vccd1 vccd1 _4986_/B sky130_fd_sc_hd__nor2_1
X_5618_ _5625_/A _5619_/B vssd1 vssd1 vccd1 vccd1 _5787_/A sky130_fd_sc_hd__nand2_2
X_6598_ _6674_/A _6634_/B vssd1 vssd1 vccd1 vccd1 _6635_/A sky130_fd_sc_hd__and2_1
X_5549_ _5581_/A _5549_/B vssd1 vssd1 vccd1 vccd1 _5551_/C sky130_fd_sc_hd__nand2_1
XFILLER_2_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7219_ _7221_/CLK hold79/X vssd1 vssd1 vccd1 vccd1 hold77/A sky130_fd_sc_hd__dfxtp_1
XFILLER_59_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_6_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7222_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_96_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4920_ _5911_/A _4913_/X _4918_/X _4919_/Y vssd1 vssd1 vccd1 vccd1 _4920_/X sky130_fd_sc_hd__a22o_1
X_4851_ _4914_/B vssd1 vssd1 vccd1 vccd1 _5880_/B sky130_fd_sc_hd__clkbuf_2
X_3802_ _4477_/A _4477_/B vssd1 vssd1 vccd1 vccd1 _3802_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4782_ _4782_/A _4782_/B vssd1 vssd1 vccd1 vccd1 _4782_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6521_ _6529_/A _6529_/B _6520_/Y vssd1 vssd1 vccd1 vccd1 _6522_/B sky130_fd_sc_hd__o21a_1
X_3733_ _3733_/A vssd1 vssd1 vccd1 vccd1 _3733_/Y sky130_fd_sc_hd__inv_2
X_3664_ _3666_/A vssd1 vssd1 vccd1 vccd1 _3664_/Y sky130_fd_sc_hd__inv_2
X_6452_ _6452_/A _6452_/B vssd1 vssd1 vccd1 vccd1 _6453_/B sky130_fd_sc_hd__and2_1
X_5403_ _5403_/A _5402_/Y vssd1 vssd1 vccd1 vccd1 _5416_/A sky130_fd_sc_hd__or2b_1
X_6383_ _6383_/A _6383_/B vssd1 vssd1 vccd1 vccd1 _6393_/B sky130_fd_sc_hd__xor2_1
X_5334_ _5213_/A _5213_/B _5216_/A vssd1 vssd1 vccd1 vccd1 _5337_/A sky130_fd_sc_hd__o21ba_1
X_5265_ _5265_/A _5265_/B vssd1 vssd1 vccd1 vccd1 _5321_/B sky130_fd_sc_hd__and2_1
X_4216_ _4216_/A _4216_/B vssd1 vssd1 vccd1 vccd1 _4218_/B sky130_fd_sc_hd__nand2_1
X_5196_ _5199_/A vssd1 vssd1 vccd1 vccd1 _6537_/B sky130_fd_sc_hd__clkbuf_2
X_7004_ _6571_/A _6993_/X _7003_/X _6995_/X vssd1 vssd1 vccd1 vccd1 _7180_/D sky130_fd_sc_hd__o211a_1
XFILLER_68_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4147_ _4147_/A _4147_/B vssd1 vssd1 vccd1 vccd1 _4149_/B sky130_fd_sc_hd__xnor2_1
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4078_ _4078_/A _4078_/B vssd1 vssd1 vccd1 vccd1 _4080_/B sky130_fd_sc_hd__nor2_1
XFILLER_24_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6719_ _6761_/B _6719_/B vssd1 vssd1 vccd1 vccd1 _6720_/B sky130_fd_sc_hd__xnor2_2
XFILLER_50_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5050_ _7175_/Q _5198_/B vssd1 vssd1 vccd1 vccd1 _5051_/A sky130_fd_sc_hd__xor2_1
X_4001_ _3910_/A _4178_/B _4000_/X vssd1 vssd1 vccd1 vccd1 _4002_/B sky130_fd_sc_hd__a21oi_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5952_ _5953_/A _5953_/B vssd1 vssd1 vccd1 vccd1 _5954_/A sky130_fd_sc_hd__nor2_1
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4903_ _4903_/A _4903_/B vssd1 vssd1 vccd1 vccd1 _4905_/A sky130_fd_sc_hd__and2_1
XFILLER_80_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5883_ _5883_/A _5883_/B vssd1 vssd1 vccd1 vccd1 _5883_/Y sky130_fd_sc_hd__nor2_1
X_4834_ _4931_/A _4931_/B _4833_/X vssd1 vssd1 vccd1 vccd1 _4837_/B sky130_fd_sc_hd__a21oi_1
XFILLER_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4765_ _7041_/A _4821_/A vssd1 vssd1 vccd1 vccd1 _4766_/B sky130_fd_sc_hd__or2_1
X_6504_ _6493_/C _5721_/A _6502_/X _6503_/X vssd1 vssd1 vccd1 vccd1 _6505_/C sky130_fd_sc_hd__a2bb2o_1
X_3716_ _3734_/A vssd1 vssd1 vccd1 vccd1 _3721_/A sky130_fd_sc_hd__buf_12
X_4696_ _4763_/A _4763_/B vssd1 vssd1 vccd1 vccd1 _4697_/B sky130_fd_sc_hd__nor2_1
X_6435_ _6483_/A _7152_/Q vssd1 vssd1 vccd1 vccd1 _6454_/B sky130_fd_sc_hd__nand2_1
X_3647_ _3647_/A vssd1 vssd1 vccd1 vccd1 _3647_/Y sky130_fd_sc_hd__inv_2
X_6366_ _6364_/X _6366_/B vssd1 vssd1 vccd1 vccd1 _6371_/A sky130_fd_sc_hd__and2b_1
XFILLER_88_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5317_ _5317_/A _5316_/A vssd1 vssd1 vccd1 vccd1 _5318_/B sky130_fd_sc_hd__or2b_1
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6297_ _6297_/A _6297_/B vssd1 vssd1 vccd1 vccd1 _6300_/A sky130_fd_sc_hd__xnor2_2
XFILLER_75_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_5248_ _5248_/A _5248_/B vssd1 vssd1 vccd1 vccd1 _5249_/B sky130_fd_sc_hd__or2_2
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold69 hold69/A vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5179_ _5325_/B _5325_/C vssd1 vssd1 vccd1 vccd1 _5180_/B sky130_fd_sc_hd__nand2_1
XFILLER_83_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4550_ _4550_/A _4550_/B vssd1 vssd1 vccd1 vccd1 _4554_/A sky130_fd_sc_hd__xor2_1
X_4481_ _4481_/A _4481_/B vssd1 vssd1 vccd1 vccd1 _4482_/B sky130_fd_sc_hd__and2_1
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6220_ _7003_/A _6329_/A _6145_/A _6145_/B vssd1 vssd1 vccd1 vccd1 _6290_/B sky130_fd_sc_hd__a22o_1
X_6151_ _7003_/A _6999_/A _6047_/B _6046_/B vssd1 vssd1 vccd1 vccd1 _6226_/B sky130_fd_sc_hd__a31o_2
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5102_ _4389_/A _4389_/B _5101_/X vssd1 vssd1 vccd1 vccd1 _5250_/B sky130_fd_sc_hd__a21oi_4
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ _6183_/A _6183_/B vssd1 vssd1 vccd1 vccd1 _6091_/A sky130_fd_sc_hd__xor2_4
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _5156_/A _5033_/B vssd1 vssd1 vccd1 vccd1 _5035_/C sky130_fd_sc_hd__xnor2_2
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6984_ _6962_/A _6977_/X _6983_/Y _6979_/X vssd1 vssd1 vccd1 vccd1 _7173_/D sky130_fd_sc_hd__o211a_1
X_5935_ _5935_/A _5935_/B vssd1 vssd1 vccd1 vccd1 _5935_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_15_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5866_ _5866_/A _5900_/A vssd1 vssd1 vccd1 vccd1 _5867_/B sky130_fd_sc_hd__or2_1
X_4817_ _4817_/A _4817_/B vssd1 vssd1 vccd1 vccd1 _4827_/A sky130_fd_sc_hd__nor2_1
X_5797_ _5798_/A _5798_/B vssd1 vssd1 vccd1 vccd1 _6076_/B sky130_fd_sc_hd__nor2_1
X_4748_ _4748_/A _4791_/A vssd1 vssd1 vccd1 vccd1 _4808_/A sky130_fd_sc_hd__xnor2_1
X_4679_ hold70/A _6627_/A vssd1 vssd1 vccd1 vccd1 _4679_/Y sky130_fd_sc_hd__nor2_1
X_6418_ _6665_/A _6691_/A _6417_/Y vssd1 vssd1 vccd1 vccd1 _6423_/A sky130_fd_sc_hd__a21o_1
X_7398_ _7398_/A _3691_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[2] sky130_fd_sc_hd__ebufn_8
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6349_ _6300_/A _6349_/B vssd1 vssd1 vccd1 vccd1 _6351_/A sky130_fd_sc_hd__and2b_1
XFILLER_88_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3981_ _5000_/B _3981_/B vssd1 vssd1 vccd1 vccd1 _5001_/B sky130_fd_sc_hd__xnor2_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5720_ _6483_/B _6439_/B vssd1 vssd1 vccd1 vccd1 _5721_/B sky130_fd_sc_hd__or2_1
XFILLER_22_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5651_ _6020_/A _5651_/B vssd1 vssd1 vccd1 vccd1 _6014_/A sky130_fd_sc_hd__nand2_1
XFILLER_30_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4602_ _4560_/B _4602_/B vssd1 vssd1 vccd1 vccd1 _4603_/B sky130_fd_sc_hd__and2b_1
X_5582_ _5557_/A _5578_/X _5581_/Y vssd1 vssd1 vccd1 vccd1 _5582_/Y sky130_fd_sc_hd__o21ai_1
X_4533_ _4533_/A _4821_/A vssd1 vssd1 vccd1 vccd1 _4766_/A sky130_fd_sc_hd__nand2_1
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4464_ _7001_/A _5812_/A vssd1 vssd1 vccd1 vccd1 _4468_/A sky130_fd_sc_hd__nor2_1
X_6203_ _6434_/B _6943_/A _6266_/B vssd1 vssd1 vccd1 vccd1 _6204_/B sky130_fd_sc_hd__mux2_2
X_4395_ _4504_/A _4504_/B _4397_/B vssd1 vssd1 vccd1 vccd1 _4407_/A sky130_fd_sc_hd__nor3_1
X_7183_ _7183_/CLK _7183_/D vssd1 vssd1 vccd1 vccd1 _7183_/Q sky130_fd_sc_hd__dfxtp_1
X_6134_ _6132_/Y _6038_/B _6133_/X vssd1 vssd1 vccd1 vccd1 _6217_/B sky130_fd_sc_hd__o21ba_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6065_ _6065_/A _5789_/A vssd1 vssd1 vccd1 vccd1 _6070_/B sky130_fd_sc_hd__or2b_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5016_ _5016_/A vssd1 vssd1 vccd1 vccd1 _7114_/A sky130_fd_sc_hd__clkbuf_2
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6967_ _7007_/A vssd1 vssd1 vccd1 vccd1 _6967_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5918_ _5918_/A _5918_/B vssd1 vssd1 vccd1 vccd1 _5950_/B sky130_fd_sc_hd__xnor2_1
XFILLER_53_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6898_ hold21/X _6892_/X _6894_/X hold41/A vssd1 vssd1 vccd1 vccd1 _6898_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5849_ _5816_/B _5849_/B vssd1 vssd1 vccd1 vccd1 _5859_/A sky130_fd_sc_hd__and2b_1
XFILLER_5_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4180_ _4694_/A _7192_/Q vssd1 vssd1 vccd1 vccd1 _4180_/X sky130_fd_sc_hd__and2_1
XFILLER_79_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6821_ _6821_/A _6821_/B vssd1 vssd1 vccd1 vccd1 _6851_/B sky130_fd_sc_hd__xnor2_2
XFILLER_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3964_ _4024_/A _4024_/B _3963_/X vssd1 vssd1 vccd1 vccd1 _3982_/A sky130_fd_sc_hd__o21a_1
X_6752_ _6750_/A _6750_/B _6750_/C vssd1 vssd1 vccd1 vccd1 _6752_/Y sky130_fd_sc_hd__a21oi_2
X_3895_ _4003_/A _7198_/Q vssd1 vssd1 vccd1 vccd1 _3896_/B sky130_fd_sc_hd__or2_1
X_6683_ _6682_/A _6681_/A _6690_/A _6665_/A vssd1 vssd1 vccd1 vccd1 _6684_/B sky130_fd_sc_hd__a22o_1
XFILLER_31_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5703_ _6049_/A _6049_/B vssd1 vssd1 vccd1 vccd1 _5710_/A sky130_fd_sc_hd__xor2_4
X_5634_ _5634_/A _5634_/B vssd1 vssd1 vccd1 vccd1 _5866_/A sky130_fd_sc_hd__xnor2_1
Xhold100 _7197_/Q vssd1 vssd1 vccd1 vccd1 _3815_/A sky130_fd_sc_hd__clkdlybuf4s50_1
X_5565_ _5575_/A _5575_/B vssd1 vssd1 vccd1 vccd1 _5567_/A sky130_fd_sc_hd__xnor2_1
X_4516_ _4516_/A _4517_/B vssd1 vssd1 vccd1 vccd1 _4601_/B sky130_fd_sc_hd__xnor2_1
Xhold111 _7016_/A vssd1 vssd1 vccd1 vccd1 hold111/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold122 hold53/X vssd1 vssd1 vccd1 vccd1 hold122/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5496_ _5496_/A _5496_/B vssd1 vssd1 vccd1 vccd1 _5497_/B sky130_fd_sc_hd__and2_1
X_4447_ _6691_/A _5854_/A vssd1 vssd1 vccd1 vccd1 _4453_/A sky130_fd_sc_hd__xnor2_2
X_7166_ _7172_/CLK _7166_/D vssd1 vssd1 vccd1 vccd1 _7166_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_98_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6117_ _6118_/B _6117_/B vssd1 vssd1 vccd1 vccd1 _6124_/C sky130_fd_sc_hd__and2_1
X_4378_ _4115_/A _4230_/A _4377_/Y vssd1 vssd1 vccd1 vccd1 _4379_/B sky130_fd_sc_hd__o21a_1
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7097_ hold82/X _7088_/X _7096_/X _7086_/X vssd1 vssd1 vccd1 vccd1 _7215_/D sky130_fd_sc_hd__o211a_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6048_ _6048_/A _6148_/B vssd1 vssd1 vccd1 vccd1 _6154_/A sky130_fd_sc_hd__xor2_4
XFILLER_73_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3680_ _3684_/A vssd1 vssd1 vccd1 vccd1 _3680_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5350_ _5350_/A _5350_/B vssd1 vssd1 vccd1 vccd1 _5351_/B sky130_fd_sc_hd__or2_1
X_5281_ _5281_/A _5394_/B vssd1 vssd1 vccd1 vccd1 _5384_/B sky130_fd_sc_hd__and2_1
X_4301_ _4301_/A _4301_/B vssd1 vssd1 vccd1 vccd1 _4370_/B sky130_fd_sc_hd__xor2_2
X_7020_ _7020_/A vssd1 vssd1 vccd1 vccd1 _7073_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4232_ _5750_/B _4232_/B vssd1 vssd1 vccd1 vccd1 _4233_/B sky130_fd_sc_hd__xor2_4
XFILLER_4_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4163_ _4163_/A _4163_/B vssd1 vssd1 vccd1 vccd1 _4164_/B sky130_fd_sc_hd__nor2_2
XFILLER_95_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4094_ _5026_/A _4573_/A _6613_/A vssd1 vssd1 vccd1 vccd1 _4094_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_67_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4996_ _3933_/A _4996_/B vssd1 vssd1 vccd1 vccd1 _4996_/X sky130_fd_sc_hd__and2b_1
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6804_ _6829_/A _6829_/B vssd1 vssd1 vccd1 vccd1 _6805_/B sky130_fd_sc_hd__xnor2_1
X_3947_ _4189_/A _4004_/A vssd1 vssd1 vccd1 vccd1 _3947_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6735_ _6763_/A _6763_/B vssd1 vssd1 vccd1 vccd1 _6736_/B sky130_fd_sc_hd__xor2_2
XFILLER_51_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6666_ _6664_/A _6664_/B _6675_/A vssd1 vssd1 vccd1 vccd1 _6667_/B sky130_fd_sc_hd__o21a_1
X_3878_ _7214_/Q vssd1 vssd1 vccd1 vccd1 _7093_/A sky130_fd_sc_hd__inv_2
X_6597_ _6597_/A _6597_/B vssd1 vssd1 vccd1 vccd1 _6634_/B sky130_fd_sc_hd__xor2_1
X_5617_ _5617_/A _5617_/B vssd1 vssd1 vccd1 vccd1 _5756_/A sky130_fd_sc_hd__nand2_4
X_5548_ _5547_/A _5547_/B _5547_/C vssd1 vssd1 vccd1 vccd1 _5549_/B sky130_fd_sc_hd__o21ai_1
X_7218_ _7221_/CLK hold73/X vssd1 vssd1 vccd1 vccd1 hold71/A sky130_fd_sc_hd__dfxtp_1
X_5479_ _5479_/A _5479_/B vssd1 vssd1 vccd1 vccd1 _5493_/A sky130_fd_sc_hd__xnor2_1
XFILLER_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7149_ _7151_/CLK hold3/X vssd1 vssd1 vccd1 vccd1 _7388_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_86_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4850_ _5913_/A vssd1 vssd1 vccd1 vccd1 _6999_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3801_ _3801_/A _3801_/B vssd1 vssd1 vccd1 vccd1 _4477_/B sky130_fd_sc_hd__xnor2_1
X_4781_ _4782_/A _4782_/B vssd1 vssd1 vccd1 vccd1 _4788_/B sky130_fd_sc_hd__xor2_1
X_6520_ _6520_/A _6520_/B vssd1 vssd1 vccd1 vccd1 _6520_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3732_ _3733_/A vssd1 vssd1 vccd1 vccd1 _3732_/Y sky130_fd_sc_hd__inv_2
X_6451_ _6452_/A _6452_/B vssd1 vssd1 vccd1 vccd1 _6453_/A sky130_fd_sc_hd__nor2_1
X_3663_ _3666_/A vssd1 vssd1 vccd1 vccd1 _3663_/Y sky130_fd_sc_hd__inv_2
X_6382_ _6395_/A _6395_/B vssd1 vssd1 vccd1 vccd1 _6383_/B sky130_fd_sc_hd__xor2_1
X_5402_ _5402_/A _5402_/B vssd1 vssd1 vccd1 vccd1 _5402_/Y sky130_fd_sc_hd__nand2_1
X_5333_ _5333_/A _5333_/B vssd1 vssd1 vccd1 vccd1 _5423_/A sky130_fd_sc_hd__xnor2_4
X_5264_ _5264_/A _5222_/A vssd1 vssd1 vccd1 vccd1 _5371_/A sky130_fd_sc_hd__or2b_1
XFILLER_87_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4215_ _4215_/A _4215_/B vssd1 vssd1 vccd1 vccd1 _4216_/B sky130_fd_sc_hd__or2_1
X_5195_ _6546_/A _5198_/B vssd1 vssd1 vccd1 vccd1 _5199_/A sky130_fd_sc_hd__nand2_1
X_7003_ _7003_/A _7011_/B vssd1 vssd1 vccd1 vccd1 _7003_/X sky130_fd_sc_hd__or2_1
XFILLER_68_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4146_ _5002_/A _4094_/Y _4092_/Y _5991_/A vssd1 vssd1 vccd1 vccd1 _4147_/B sky130_fd_sc_hd__o2bb2a_2
XFILLER_95_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4077_ _4054_/A _4053_/B _4070_/A vssd1 vssd1 vccd1 vccd1 _4078_/B sky130_fd_sc_hd__o21ba_1
XFILLER_36_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4979_ _4979_/A _4979_/B vssd1 vssd1 vccd1 vccd1 _4995_/A sky130_fd_sc_hd__nor2_1
X_6718_ _6718_/A _6718_/B vssd1 vssd1 vccd1 vccd1 _6778_/B sky130_fd_sc_hd__nor2_1
X_6649_ _6649_/A _6649_/B vssd1 vssd1 vccd1 vccd1 _6706_/B sky130_fd_sc_hd__nor2_1
XFILLER_50_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4000_ _4392_/B _7194_/Q vssd1 vssd1 vccd1 vccd1 _4000_/X sky130_fd_sc_hd__and2_1
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5951_ _5955_/B _5955_/A vssd1 vssd1 vccd1 vccd1 _5957_/A sky130_fd_sc_hd__or2b_1
XFILLER_65_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4902_ _4902_/A _4902_/B vssd1 vssd1 vccd1 vccd1 _4903_/B sky130_fd_sc_hd__or2_1
X_5882_ _5883_/A _5883_/B vssd1 vssd1 vccd1 vccd1 _5908_/B sky130_fd_sc_hd__xor2_1
XFILLER_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4833_ _4832_/B _4833_/B vssd1 vssd1 vccd1 vccd1 _4833_/X sky130_fd_sc_hd__and2b_1
XFILLER_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4764_ _4822_/B _4768_/C vssd1 vssd1 vccd1 vccd1 _4820_/A sky130_fd_sc_hd__xnor2_2
X_6503_ _6502_/B _5691_/B _6484_/B vssd1 vssd1 vccd1 vccd1 _6503_/X sky130_fd_sc_hd__a21o_1
X_3715_ _3715_/A vssd1 vssd1 vccd1 vccd1 _3715_/Y sky130_fd_sc_hd__inv_2
X_4695_ _4695_/A _4695_/B vssd1 vssd1 vccd1 vccd1 _4761_/A sky130_fd_sc_hd__xor2_2
X_6434_ _6434_/A _6434_/B vssd1 vssd1 vccd1 vccd1 _6454_/A sky130_fd_sc_hd__xnor2_1
X_3646_ _3647_/A vssd1 vssd1 vccd1 vccd1 _3646_/Y sky130_fd_sc_hd__inv_2
X_6365_ _6365_/A _6365_/B _6363_/X vssd1 vssd1 vccd1 vccd1 _6366_/B sky130_fd_sc_hd__or3b_1
X_6296_ _6296_/A vssd1 vssd1 vccd1 vccd1 _6297_/B sky130_fd_sc_hd__inv_2
X_5316_ _5316_/A _5317_/A vssd1 vssd1 vccd1 vccd1 _5318_/A sky130_fd_sc_hd__or2b_1
X_5247_ _5095_/A _5247_/B vssd1 vssd1 vccd1 vccd1 _5248_/B sky130_fd_sc_hd__and2b_1
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_5178_ _5178_/A _5178_/B vssd1 vssd1 vccd1 vccd1 _5325_/C sky130_fd_sc_hd__nand2_1
XFILLER_28_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4129_ _7167_/Q _5688_/A vssd1 vssd1 vccd1 vccd1 _4133_/A sky130_fd_sc_hd__or2_1
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4480_ _5625_/A vssd1 vssd1 vccd1 vccd1 _6624_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6150_ _6223_/B _6150_/B vssd1 vssd1 vccd1 vccd1 _6153_/A sky130_fd_sc_hd__xnor2_4
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _4390_/B _5101_/B vssd1 vssd1 vccd1 vccd1 _5101_/X sky130_fd_sc_hd__and2b_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ _5811_/A _5811_/B _6080_/X vssd1 vssd1 vccd1 vccd1 _6183_/B sky130_fd_sc_hd__a21oi_4
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _5032_/A _5032_/B vssd1 vssd1 vccd1 vccd1 _5033_/B sky130_fd_sc_hd__xor2_1
XFILLER_65_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6983_ _6983_/A _6983_/B vssd1 vssd1 vccd1 vccd1 _6983_/Y sky130_fd_sc_hd__nand2_1
XFILLER_15_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5934_ _5934_/A _6100_/B vssd1 vssd1 vccd1 vccd1 _6011_/A sky130_fd_sc_hd__xnor2_1
X_5865_ _5865_/A _5865_/B vssd1 vssd1 vccd1 vccd1 _5890_/A sky130_fd_sc_hd__xnor2_1
X_4816_ _4816_/A _4816_/B vssd1 vssd1 vccd1 vccd1 _4817_/B sky130_fd_sc_hd__and2_1
X_5796_ _6805_/A _5796_/B vssd1 vssd1 vccd1 vccd1 _5798_/B sky130_fd_sc_hd__xor2_1
X_4747_ _4790_/A _4790_/B vssd1 vssd1 vccd1 vccd1 _4791_/A sky130_fd_sc_hd__nor2_1
X_4678_ _4684_/A _4678_/B vssd1 vssd1 vccd1 vccd1 _4739_/A sky130_fd_sc_hd__xnor2_1
X_7397_ _7397_/A _3690_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[1] sky130_fd_sc_hd__ebufn_8
X_6417_ _6560_/A _6417_/B vssd1 vssd1 vccd1 vccd1 _6417_/Y sky130_fd_sc_hd__nor2_1
X_3629_ _3629_/A vssd1 vssd1 vccd1 vccd1 _3629_/Y sky130_fd_sc_hd__inv_2
X_6348_ _6348_/A _6348_/B vssd1 vssd1 vccd1 vccd1 _6385_/B sky130_fd_sc_hd__xnor2_1
XFILLER_76_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6279_ _6213_/A _6213_/B _6215_/A _6215_/B vssd1 vssd1 vccd1 vccd1 _6280_/B sky130_fd_sc_hd__o22a_1
XFILLER_48_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3980_ _3980_/A _3980_/B vssd1 vssd1 vccd1 vccd1 _3981_/B sky130_fd_sc_hd__xnor2_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5650_ _7157_/Q _6494_/B vssd1 vssd1 vccd1 vccd1 _5651_/B sky130_fd_sc_hd__or2b_1
X_4601_ _4601_/A _4601_/B vssd1 vssd1 vccd1 vccd1 _4625_/A sky130_fd_sc_hd__xnor2_1
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5581_ _5581_/A _5581_/B vssd1 vssd1 vccd1 vccd1 _5581_/Y sky130_fd_sc_hd__xnor2_1
X_4532_ _7192_/Q vssd1 vssd1 vccd1 vccd1 _4821_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4463_ _5872_/A vssd1 vssd1 vccd1 vccd1 _7001_/A sky130_fd_sc_hd__inv_2
X_6202_ _6464_/B vssd1 vssd1 vccd1 vccd1 _6943_/A sky130_fd_sc_hd__clkbuf_2
X_4394_ _7083_/A _4394_/B vssd1 vssd1 vccd1 vccd1 _4397_/B sky130_fd_sc_hd__xnor2_2
X_7182_ _7183_/CLK _7182_/D vssd1 vssd1 vccd1 vccd1 _7182_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6133_ _6037_/A _6133_/B vssd1 vssd1 vccd1 vccd1 _6133_/X sky130_fd_sc_hd__and2b_1
X_6064_ _6064_/A _6180_/A vssd1 vssd1 vccd1 vccd1 _6073_/A sky130_fd_sc_hd__nor2_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _5015_/A _5015_/B vssd1 vssd1 vccd1 vccd1 _5156_/A sky130_fd_sc_hd__xnor2_2
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6966_ _6966_/A _6983_/B vssd1 vssd1 vccd1 vccd1 _6966_/Y sky130_fd_sc_hd__nand2_1
X_5917_ _5948_/A _5945_/A vssd1 vssd1 vccd1 vccd1 _5918_/B sky130_fd_sc_hd__and2b_1
XFILLER_53_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6897_ _6906_/A hold39/X vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__nor2_1
X_5848_ _5643_/A _5643_/B _5647_/B vssd1 vssd1 vccd1 vccd1 _5861_/A sky130_fd_sc_hd__a21oi_4
X_5779_ _5822_/A _5777_/X _5778_/X vssd1 vssd1 vccd1 vccd1 _5780_/B sky130_fd_sc_hd__o21a_1
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7271__64 vssd1 vssd1 vccd1 vccd1 _7271__64/HI _7370_/A sky130_fd_sc_hd__conb_1
XFILLER_44_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6820_ _6112_/A _6796_/B _6799_/B _6111_/B vssd1 vssd1 vccd1 vccd1 _6821_/B sky130_fd_sc_hd__o211a_1
XFILLER_35_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3963_ _3963_/A _3963_/B vssd1 vssd1 vccd1 vccd1 _3963_/X sky130_fd_sc_hd__or2_1
X_6751_ _6751_/A vssd1 vssd1 vccd1 vccd1 _6751_/Y sky130_fd_sc_hd__inv_2
X_3894_ _4526_/B _4873_/A vssd1 vssd1 vccd1 vccd1 _3904_/A sky130_fd_sc_hd__nand2_1
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_6682_ _6682_/A _6682_/B vssd1 vssd1 vccd1 vccd1 _6690_/A sky130_fd_sc_hd__xor2_2
X_5702_ _5715_/A _5715_/B _5716_/B _5701_/Y vssd1 vssd1 vccd1 vccd1 _6049_/B sky130_fd_sc_hd__a31oi_4
X_5633_ _5634_/B _5634_/A vssd1 vssd1 vccd1 vccd1 _5863_/A sky130_fd_sc_hd__or2b_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5564_ _5564_/A _5564_/B vssd1 vssd1 vccd1 vccd1 _5575_/B sky130_fd_sc_hd__nand2_1
X_4515_ _4604_/A _4604_/B _4514_/X vssd1 vssd1 vccd1 vccd1 _4517_/B sky130_fd_sc_hd__a21o_1
Xhold101 _7071_/X vssd1 vssd1 vccd1 vccd1 _7205_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold123 _5829_/B vssd1 vssd1 vccd1 vccd1 hold123/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_5495_ _5496_/A _5496_/B vssd1 vssd1 vccd1 vccd1 _5556_/A sky130_fd_sc_hd__nor2_1
Xhold112 _5762_/A vssd1 vssd1 vccd1 vccd1 hold112/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_4446_ _4450_/B vssd1 vssd1 vccd1 vccd1 _6691_/A sky130_fd_sc_hd__buf_2
X_7165_ _7172_/CLK _7165_/D vssd1 vssd1 vccd1 vccd1 _7165_/Q sky130_fd_sc_hd__dfxtp_2
X_4377_ _6713_/A _4377_/B vssd1 vssd1 vccd1 vccd1 _4377_/Y sky130_fd_sc_hd__nand2_1
XFILLER_98_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6116_ _6128_/B _6116_/B vssd1 vssd1 vccd1 vccd1 _6124_/A sky130_fd_sc_hd__and2b_1
XFILLER_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7096_ _7096_/A _7106_/B vssd1 vssd1 vccd1 vccd1 _7096_/X sky130_fd_sc_hd__or2_1
XFILLER_58_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6047_ _6047_/A _6047_/B vssd1 vssd1 vccd1 vccd1 _6148_/B sky130_fd_sc_hd__xnor2_2
XFILLER_100_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6949_ _6977_/A vssd1 vssd1 vccd1 vccd1 _6949_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7321__114 vssd1 vssd1 vccd1 vccd1 _7321__114/HI _7429_/A sky130_fd_sc_hd__conb_1
XFILLER_1_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4300_ _4379_/A _4300_/B vssd1 vssd1 vccd1 vccd1 _4301_/B sky130_fd_sc_hd__xnor2_1
X_5280_ _7055_/A _5280_/B vssd1 vssd1 vccd1 vccd1 _5394_/B sky130_fd_sc_hd__or2_1
XFILLER_99_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4231_ _6713_/A _4296_/B vssd1 vssd1 vccd1 vccd1 _4232_/B sky130_fd_sc_hd__xnor2_4
XFILLER_67_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4162_ _4162_/A _4162_/B vssd1 vssd1 vccd1 vccd1 _4163_/B sky130_fd_sc_hd__and2_1
XFILLER_95_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4093_ _4329_/A vssd1 vssd1 vccd1 vccd1 _5026_/A sky130_fd_sc_hd__inv_2
XFILLER_48_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4995_ _4995_/A _4995_/B vssd1 vssd1 vccd1 vccd1 _4998_/A sky130_fd_sc_hd__xnor2_1
XFILLER_23_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6803_ _6981_/A _6771_/B _6802_/Y vssd1 vssd1 vccd1 vccd1 _6829_/B sky130_fd_sc_hd__o21a_1
XFILLER_51_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3946_ _4189_/A _4004_/A vssd1 vssd1 vccd1 vccd1 _4026_/B sky130_fd_sc_hd__xor2_2
X_6734_ _6852_/A _6527_/B _6733_/X vssd1 vssd1 vccd1 vccd1 _6763_/B sky130_fd_sc_hd__a21oi_2
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6665_ _6665_/A _6674_/B vssd1 vssd1 vccd1 vccd1 _6675_/A sky130_fd_sc_hd__nand2_1
X_3877_ _3879_/B _5276_/A _3877_/C vssd1 vssd1 vccd1 vccd1 _3889_/B sky130_fd_sc_hd__and3_1
X_6596_ _6736_/A _6596_/B vssd1 vssd1 vccd1 vccd1 _6597_/B sky130_fd_sc_hd__xnor2_1
X_5616_ _6983_/A _5895_/A vssd1 vssd1 vccd1 vccd1 _5617_/B sky130_fd_sc_hd__nand2_1
X_5547_ _5547_/A _5547_/B _5547_/C vssd1 vssd1 vccd1 vccd1 _5581_/A sky130_fd_sc_hd__or3_1
XFILLER_2_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5478_ _5478_/A _5541_/B vssd1 vssd1 vccd1 vccd1 _5479_/B sky130_fd_sc_hd__xnor2_2
X_7217_ _7221_/CLK _7217_/D vssd1 vssd1 vccd1 vccd1 _7217_/Q sky130_fd_sc_hd__dfxtp_1
X_4429_ _4429_/A _4429_/B vssd1 vssd1 vccd1 vccd1 _4550_/A sky130_fd_sc_hd__xnor2_2
XFILLER_58_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7148_ _7226_/CLK hold11/X vssd1 vssd1 vccd1 vccd1 _7387_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_48_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7079_ hold97/X _7075_/X _7078_/X _7073_/X vssd1 vssd1 vccd1 vccd1 _7208_/D sky130_fd_sc_hd__o211a_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7241__34 vssd1 vssd1 vccd1 vccd1 _7241__34/HI _7340_/A sky130_fd_sc_hd__conb_1
XFILLER_64_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4780_ _4812_/A _4812_/B _4779_/X vssd1 vssd1 vccd1 vccd1 _4782_/B sky130_fd_sc_hd__a21oi_1
X_3800_ _5347_/A _6120_/B vssd1 vssd1 vccd1 vccd1 _4477_/A sky130_fd_sc_hd__nand2_2
X_3731_ _3733_/A vssd1 vssd1 vccd1 vccd1 _3731_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3662_ _3666_/A vssd1 vssd1 vccd1 vccd1 _3662_/Y sky130_fd_sc_hd__inv_2
X_6450_ _6464_/B _6112_/A _6449_/Y vssd1 vssd1 vccd1 vccd1 _6452_/B sky130_fd_sc_hd__a21oi_1
XFILLER_9_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6381_ _6379_/X _6348_/B _6380_/X vssd1 vssd1 vccd1 vccd1 _6395_/B sky130_fd_sc_hd__a21oi_1
X_5401_ _5402_/A _5402_/B vssd1 vssd1 vccd1 vccd1 _5403_/A sky130_fd_sc_hd__nor2_1
X_5332_ _6539_/A _5332_/B vssd1 vssd1 vccd1 vccd1 _5333_/B sky130_fd_sc_hd__xnor2_2
X_5263_ _5263_/A _5256_/A vssd1 vssd1 vccd1 vccd1 _5375_/A sky130_fd_sc_hd__or2b_1
X_4214_ _4409_/A _4408_/B _4408_/A vssd1 vssd1 vccd1 vccd1 _4218_/A sky130_fd_sc_hd__a21boi_2
X_5194_ _7175_/Q vssd1 vssd1 vccd1 vccd1 _6802_/A sky130_fd_sc_hd__inv_2
X_7002_ _6736_/A _6993_/X _7001_/Y _6995_/X vssd1 vssd1 vccd1 vccd1 _7179_/D sky130_fd_sc_hd__o211a_1
X_4145_ _4573_/A vssd1 vssd1 vccd1 vccd1 _5991_/A sky130_fd_sc_hd__buf_2
XFILLER_83_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4076_ hold77/A _4076_/B _4076_/C vssd1 vssd1 vccd1 vccd1 _4197_/A sky130_fd_sc_hd__nor3_1
XFILLER_83_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4978_ _4978_/A _4978_/B _4978_/C vssd1 vssd1 vccd1 vccd1 _4979_/B sky130_fd_sc_hd__and3_1
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3929_ _4008_/A _4008_/B _3928_/X vssd1 vssd1 vccd1 vccd1 _3931_/B sky130_fd_sc_hd__a21o_1
X_6717_ _6717_/A _6717_/B vssd1 vssd1 vccd1 vccd1 _6778_/A sky130_fd_sc_hd__nor2_1
X_6648_ _6649_/A _6649_/B vssd1 vssd1 vccd1 vccd1 _6706_/A sky130_fd_sc_hd__and2_1
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6579_ _6579_/A _6579_/B vssd1 vssd1 vccd1 vccd1 _6580_/B sky130_fd_sc_hd__xnor2_1
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5950_ _5950_/A _5950_/B vssd1 vssd1 vccd1 vccd1 _5955_/A sky130_fd_sc_hd__xnor2_1
X_4901_ _4904_/A _4904_/B vssd1 vssd1 vccd1 vccd1 _4906_/A sky130_fd_sc_hd__and2b_1
XFILLER_80_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5881_ _5879_/A _5878_/Y _5910_/A vssd1 vssd1 vccd1 vccd1 _5883_/B sky130_fd_sc_hd__a21oi_2
X_4832_ _4833_/B _4832_/B vssd1 vssd1 vccd1 vccd1 _4931_/B sky130_fd_sc_hd__xnor2_1
X_4763_ _4763_/A _4763_/B vssd1 vssd1 vccd1 vccd1 _4768_/C sky130_fd_sc_hd__xor2_2
XFILLER_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4694_ _4694_/A _4694_/B vssd1 vssd1 vccd1 vccd1 _4763_/B sky130_fd_sc_hd__xnor2_2
X_6502_ _6502_/A _6502_/B vssd1 vssd1 vccd1 vccd1 _6502_/X sky130_fd_sc_hd__xor2_1
X_3714_ _3715_/A vssd1 vssd1 vccd1 vccd1 _3714_/Y sky130_fd_sc_hd__inv_2
X_6433_ _4429_/A _4553_/A _6588_/A _6441_/C vssd1 vssd1 vccd1 vccd1 _6481_/A sky130_fd_sc_hd__a31o_1
X_3645_ _3647_/A vssd1 vssd1 vccd1 vccd1 _3645_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6364_ _6365_/A _6365_/B _6363_/X vssd1 vssd1 vccd1 vccd1 _6364_/X sky130_fd_sc_hd__o21ba_1
XFILLER_88_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6295_ _6295_/A _6346_/C vssd1 vssd1 vccd1 vccd1 _6296_/A sky130_fd_sc_hd__or2_1
X_5315_ _5315_/A _5315_/B vssd1 vssd1 vccd1 vccd1 _5317_/A sky130_fd_sc_hd__xnor2_1
XFILLER_88_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5246_ _5094_/B _5246_/B vssd1 vssd1 vccd1 vccd1 _5248_/A sky130_fd_sc_hd__and2b_1
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_28_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5177_ _5178_/A _5178_/B vssd1 vssd1 vccd1 vccd1 _5325_/B sky130_fd_sc_hd__or2_1
XFILLER_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4128_ _4286_/A _6039_/B vssd1 vssd1 vccd1 vccd1 _5688_/A sky130_fd_sc_hd__and2_2
X_4059_ _4794_/A vssd1 vssd1 vccd1 vccd1 _5597_/B sky130_fd_sc_hd__buf_2
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6080_ _5780_/B _6080_/B vssd1 vssd1 vccd1 vccd1 _6080_/X sky130_fd_sc_hd__and2b_1
X_5100_ _5100_/A _5100_/B vssd1 vssd1 vccd1 vccd1 _5250_/A sky130_fd_sc_hd__xnor2_2
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _4159_/A _4158_/B _4158_/A vssd1 vssd1 vccd1 vccd1 _5032_/B sky130_fd_sc_hd__o21ba_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7277__70 vssd1 vssd1 vccd1 vccd1 _7277__70/HI _7376_/A sky130_fd_sc_hd__conb_1
XFILLER_85_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6982_ _6960_/A _6977_/X _6981_/Y _6979_/X vssd1 vssd1 vccd1 vccd1 _7172_/D sky130_fd_sc_hd__o211a_1
XFILLER_53_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5933_ _5930_/A _5930_/B _5935_/B _5935_/A vssd1 vssd1 vccd1 vccd1 _6100_/B sky130_fd_sc_hd__a2bb2o_2
X_5864_ _5893_/A _5864_/B vssd1 vssd1 vccd1 vccd1 _5894_/A sky130_fd_sc_hd__nor2_1
X_4815_ _4815_/A _4815_/B vssd1 vssd1 vccd1 vccd1 _4869_/A sky130_fd_sc_hd__xnor2_1
XFILLER_31_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5795_ _6850_/A _5795_/B vssd1 vssd1 vccd1 vccd1 _6805_/A sky130_fd_sc_hd__nand2_4
X_4746_ _6137_/B _4746_/B vssd1 vssd1 vccd1 vccd1 _4790_/B sky130_fd_sc_hd__xnor2_1
X_4677_ _4672_/Y _4742_/B _4676_/Y vssd1 vssd1 vccd1 vccd1 _4678_/B sky130_fd_sc_hd__o21a_1
X_3628_ _3629_/A vssd1 vssd1 vccd1 vccd1 _3628_/Y sky130_fd_sc_hd__inv_2
X_6416_ _5936_/A _4330_/A _4328_/B vssd1 vssd1 vccd1 vccd1 _6417_/B sky130_fd_sc_hd__o21ai_2
X_7396_ _7396_/A _3735_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[0] sky130_fd_sc_hd__ebufn_8
X_6347_ _6383_/A _6347_/B vssd1 vssd1 vccd1 vccd1 _6348_/B sky130_fd_sc_hd__nor2_1
XFILLER_88_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6278_ _6325_/A _6325_/B vssd1 vssd1 vccd1 vccd1 _6280_/A sky130_fd_sc_hd__xnor2_2
X_5229_ _5229_/A _5229_/B _5229_/C vssd1 vssd1 vccd1 vccd1 _5231_/A sky130_fd_sc_hd__and3_1
XFILLER_84_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_94_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4600_ _4600_/A _4600_/B vssd1 vssd1 vccd1 vccd1 _4688_/A sky130_fd_sc_hd__xor2_1
X_5580_ _7011_/A _5486_/Y _5542_/A vssd1 vssd1 vccd1 vccd1 _5581_/B sky130_fd_sc_hd__o21ba_1
X_4531_ _7043_/A _4531_/B vssd1 vssd1 vccd1 vccd1 _4535_/A sky130_fd_sc_hd__xnor2_1
X_4462_ _4466_/A vssd1 vssd1 vccd1 vccd1 _5872_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6201_ _7158_/Q _7157_/Q vssd1 vssd1 vccd1 vccd1 _6434_/B sky130_fd_sc_hd__xor2_2
XFILLER_98_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4393_ _4393_/A _4393_/B vssd1 vssd1 vccd1 vccd1 _4504_/B sky130_fd_sc_hd__nand2_1
X_7181_ _7183_/CLK _7181_/D vssd1 vssd1 vccd1 vccd1 _7181_/Q sky130_fd_sc_hd__dfxtp_1
X_6132_ _6132_/A vssd1 vssd1 vccd1 vccd1 _6132_/Y sky130_fd_sc_hd__inv_2
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6063_ _6063_/A _6063_/B _6063_/C vssd1 vssd1 vccd1 vccd1 _6180_/A sky130_fd_sc_hd__nor3_1
X_5014_ _5228_/B _5014_/B vssd1 vssd1 vccd1 vccd1 _5015_/B sky130_fd_sc_hd__xor2_2
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6965_ _7080_/A vssd1 vssd1 vccd1 vccd1 _6983_/B sky130_fd_sc_hd__buf_2
XFILLER_53_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5916_ _6994_/A _5944_/B vssd1 vssd1 vccd1 vccd1 _5945_/A sky130_fd_sc_hd__nor2_1
XFILLER_34_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6896_ hold28/X _6890_/X _6895_/X vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__a21oi_1
XFILLER_22_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5847_ _6092_/A _6092_/B vssd1 vssd1 vccd1 vccd1 _5862_/A sky130_fd_sc_hd__xor2_2
X_5778_ _5821_/A _5821_/B vssd1 vssd1 vccd1 vccd1 _5778_/X sky130_fd_sc_hd__or2_1
X_4729_ _4802_/A vssd1 vssd1 vccd1 vccd1 _4770_/A sky130_fd_sc_hd__inv_2
XFILLER_89_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7379_ _7379_/A _3669_/Y vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__ebufn_8
XFILLER_88_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7247__40 vssd1 vssd1 vccd1 vccd1 _7247__40/HI _7346_/A sky130_fd_sc_hd__conb_1
XFILLER_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6750_ _6750_/A _6750_/B _6750_/C vssd1 vssd1 vccd1 vccd1 _6751_/A sky130_fd_sc_hd__nand3_2
XFILLER_23_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3962_ _4157_/B _3962_/B vssd1 vssd1 vccd1 vccd1 _4024_/B sky130_fd_sc_hd__nand2_2
X_5701_ _5698_/A _5698_/B _5700_/B vssd1 vssd1 vccd1 vccd1 _5701_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_50_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3893_ _7184_/Q vssd1 vssd1 vccd1 vccd1 _4873_/A sky130_fd_sc_hd__clkbuf_2
X_6681_ _6681_/A _6577_/A vssd1 vssd1 vccd1 vccd1 _6682_/B sky130_fd_sc_hd__or2b_1
XFILLER_31_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5632_ _5630_/A _5812_/B _5631_/X vssd1 vssd1 vccd1 vccd1 _5634_/A sky130_fd_sc_hd__a21bo_1
X_5563_ _5563_/A _5563_/B vssd1 vssd1 vccd1 vccd1 _5564_/B sky130_fd_sc_hd__nand2_1
X_4514_ _4514_/A _4514_/B vssd1 vssd1 vccd1 vccd1 _4514_/X sky130_fd_sc_hd__and2_1
Xhold124 _4412_/A vssd1 vssd1 vccd1 vccd1 hold124/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold113 _6479_/B vssd1 vssd1 vccd1 vccd1 _6929_/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold102 _4527_/A vssd1 vssd1 vccd1 vccd1 _4400_/A sky130_fd_sc_hd__clkbuf_2
X_5494_ _5402_/Y _5416_/B _5403_/A vssd1 vssd1 vccd1 vccd1 _5496_/B sky130_fd_sc_hd__a21oi_1
X_4445_ _4445_/A _4445_/B vssd1 vssd1 vccd1 vccd1 _4488_/A sky130_fd_sc_hd__xnor2_1
X_7164_ _7172_/CLK _7164_/D vssd1 vssd1 vccd1 vccd1 _7164_/Q sky130_fd_sc_hd__dfxtp_1
X_4376_ _5229_/A _4375_/Y _4298_/Y vssd1 vssd1 vccd1 vccd1 _4380_/A sky130_fd_sc_hd__o21ai_1
XFILLER_100_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6115_ _6115_/A _6115_/B vssd1 vssd1 vccd1 vccd1 _6210_/A sky130_fd_sc_hd__xor2_4
XFILLER_58_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7095_ _7095_/A vssd1 vssd1 vccd1 vccd1 _7106_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6046_ _6046_/A _6046_/B vssd1 vssd1 vccd1 vccd1 _6047_/B sky130_fd_sc_hd__nor2_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6948_ _6926_/A _6935_/X _6947_/Y _6939_/X vssd1 vssd1 vccd1 vccd1 _7160_/D sky130_fd_sc_hd__o211a_1
X_6879_ _6879_/A hold65/A vssd1 vssd1 vccd1 vccd1 hold64/A sky130_fd_sc_hd__nand2_1
XFILLER_22_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4230_ _4230_/A _4230_/B vssd1 vssd1 vccd1 vccd1 _4296_/B sky130_fd_sc_hd__and2_1
X_4161_ _4162_/A _4162_/B vssd1 vssd1 vccd1 vccd1 _4163_/A sky130_fd_sc_hd__nor2_1
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4092_ _5019_/A _6613_/A vssd1 vssd1 vccd1 vccd1 _4092_/Y sky130_fd_sc_hd__nand2_2
XFILLER_82_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6802_ _6802_/A _6802_/B vssd1 vssd1 vccd1 vccd1 _6802_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4994_ _4994_/A _4994_/B vssd1 vssd1 vccd1 vccd1 _4995_/B sky130_fd_sc_hd__xor2_1
X_3945_ _7208_/Q _4003_/A vssd1 vssd1 vccd1 vccd1 _4004_/A sky130_fd_sc_hd__or2b_2
X_6733_ _6526_/A _6733_/B vssd1 vssd1 vccd1 vccd1 _6733_/X sky130_fd_sc_hd__and2b_1
XFILLER_51_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6664_ _6664_/A _6664_/B vssd1 vssd1 vccd1 vccd1 _6674_/B sky130_fd_sc_hd__xor2_1
X_3876_ _4957_/A vssd1 vssd1 vccd1 vccd1 _5276_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5615_ _5615_/A vssd1 vssd1 vccd1 vccd1 _6983_/A sky130_fd_sc_hd__clkbuf_4
X_6595_ _6620_/A _6620_/B _6594_/X vssd1 vssd1 vccd1 vccd1 _6597_/A sky130_fd_sc_hd__a21oi_1
X_5546_ _5546_/A _5492_/B vssd1 vssd1 vccd1 vccd1 _5551_/B sky130_fd_sc_hd__or2b_1
XFILLER_2_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5477_ _5399_/A _5399_/B _5387_/A vssd1 vssd1 vccd1 vccd1 _5479_/A sky130_fd_sc_hd__a21oi_2
X_4428_ _4208_/A _6479_/B _4641_/A vssd1 vssd1 vccd1 vccd1 _4429_/B sky130_fd_sc_hd__a21oi_1
X_7216_ _7221_/CLK _7216_/D vssd1 vssd1 vccd1 vccd1 hold80/A sky130_fd_sc_hd__dfxtp_1
XFILLER_86_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4359_ _4359_/A _4359_/B vssd1 vssd1 vccd1 vccd1 _5057_/B sky130_fd_sc_hd__or2_1
X_7147_ _7151_/CLK _7147_/D vssd1 vssd1 vccd1 vccd1 _7386_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7078_ _7078_/A _7091_/B vssd1 vssd1 vccd1 vccd1 _7078_/X sky130_fd_sc_hd__or2_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6029_ _6029_/A _6029_/B vssd1 vssd1 vccd1 vccd1 _6117_/B sky130_fd_sc_hd__nor2_1
XFILLER_39_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3730_ _3733_/A vssd1 vssd1 vccd1 vccd1 _3730_/Y sky130_fd_sc_hd__inv_2
X_3661_ _3679_/A vssd1 vssd1 vccd1 vccd1 _3666_/A sky130_fd_sc_hd__buf_12
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6380_ _6344_/A _6380_/B vssd1 vssd1 vccd1 vccd1 _6380_/X sky130_fd_sc_hd__and2b_1
X_5400_ _5295_/A _5295_/B _5285_/A vssd1 vssd1 vccd1 vccd1 _5402_/B sky130_fd_sc_hd__a21oi_1
X_5331_ _5202_/A _5330_/Y _5200_/Y vssd1 vssd1 vccd1 vccd1 _5332_/B sky130_fd_sc_hd__a21oi_1
X_5262_ _6261_/A vssd1 vssd1 vccd1 vccd1 _5262_/X sky130_fd_sc_hd__clkbuf_2
X_7001_ _7001_/A _7006_/B vssd1 vssd1 vccd1 vccd1 _7001_/Y sky130_fd_sc_hd__nand2_1
X_4213_ _7089_/A hold71/A _7217_/Q vssd1 vssd1 vccd1 vccd1 _4408_/A sky130_fd_sc_hd__or3_1
X_5193_ _7175_/Q _6564_/A _6546_/A vssd1 vssd1 vccd1 vccd1 _5193_/X sky130_fd_sc_hd__a21o_1
XFILLER_95_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4144_ _4139_/Y _6063_/B _4143_/X vssd1 vssd1 vccd1 vccd1 _4147_/A sky130_fd_sc_hd__a21o_1
XFILLER_95_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4075_ hold96/A _4721_/A vssd1 vssd1 vccd1 vccd1 _4076_/C sky130_fd_sc_hd__nor2_1
XFILLER_70_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4977_ _4978_/A _4978_/B _4978_/C vssd1 vssd1 vccd1 vccd1 _4979_/A sky130_fd_sc_hd__a21oi_1
X_6716_ _6793_/A _6716_/B vssd1 vssd1 vccd1 vccd1 _6744_/A sky130_fd_sc_hd__or2_1
X_3928_ _3927_/B _3928_/B vssd1 vssd1 vccd1 vccd1 _3928_/X sky130_fd_sc_hd__and2b_1
X_3859_ _4950_/A _4950_/B vssd1 vssd1 vccd1 vccd1 _4951_/A sky130_fd_sc_hd__xor2_1
X_6647_ _6647_/A _6647_/B vssd1 vssd1 vccd1 vccd1 _6707_/A sky130_fd_sc_hd__xnor2_2
XFILLER_50_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6578_ _6576_/A _6576_/B _6603_/A vssd1 vssd1 vccd1 vccd1 _6581_/B sky130_fd_sc_hd__a21o_1
XFILLER_3_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5529_ _5529_/A _5529_/B vssd1 vssd1 vccd1 vccd1 _5530_/B sky130_fd_sc_hd__nand2_1
XFILLER_1_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7301__94 vssd1 vssd1 vccd1 vccd1 _7301__94/HI _7409_/A sky130_fd_sc_hd__conb_1
XFILLER_101_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4900_ _4917_/B _4919_/B _4899_/Y vssd1 vssd1 vccd1 vccd1 _4904_/B sky130_fd_sc_hd__a21o_1
XFILLER_80_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5880_ _5824_/A _5880_/B _5880_/C vssd1 vssd1 vccd1 vccd1 _5910_/A sky130_fd_sc_hd__and3b_1
XFILLER_65_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4831_ _4928_/A _4927_/B _4927_/A vssd1 vssd1 vccd1 vccd1 _4832_/B sky130_fd_sc_hd__o21ba_1
XFILLER_33_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4762_ _4821_/A _4821_/B vssd1 vssd1 vccd1 vccd1 _4822_/B sky130_fd_sc_hd__nand2_2
X_3713_ _3715_/A vssd1 vssd1 vccd1 vccd1 _3713_/Y sky130_fd_sc_hd__inv_2
X_6501_ _6496_/A _6496_/C _6496_/B vssd1 vssd1 vccd1 vccd1 _6505_/B sky130_fd_sc_hd__o21ai_1
X_4693_ _4693_/A _4693_/B vssd1 vssd1 vccd1 vccd1 _4697_/A sky130_fd_sc_hd__xnor2_2
X_6432_ _6445_/B _6432_/B _6432_/C vssd1 vssd1 vccd1 vccd1 _6441_/C sky130_fd_sc_hd__and3_1
X_3644_ _3647_/A vssd1 vssd1 vccd1 vccd1 _3644_/Y sky130_fd_sc_hd__inv_2
X_6363_ _6327_/A _6327_/B _6330_/A _6270_/X vssd1 vssd1 vccd1 vccd1 _6363_/X sky130_fd_sc_hd__o211a_1
X_6294_ _6293_/B _6294_/B vssd1 vssd1 vccd1 vccd1 _6346_/C sky130_fd_sc_hd__and2b_1
X_5314_ _5314_/A _5314_/B vssd1 vssd1 vccd1 vccd1 _5315_/B sky130_fd_sc_hd__xnor2_2
XFILLER_29_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5245_ _5245_/A _5368_/B vssd1 vssd1 vccd1 vccd1 _5249_/A sky130_fd_sc_hd__xnor2_4
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_5176_ _5176_/A _5176_/B vssd1 vssd1 vccd1 vccd1 _5178_/B sky130_fd_sc_hd__xor2_1
XFILLER_83_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4127_ _4374_/A _5011_/A vssd1 vssd1 vccd1 vccd1 _6039_/B sky130_fd_sc_hd__or2_1
X_4058_ _4794_/A _6449_/A vssd1 vssd1 vccd1 vccd1 _5017_/A sky130_fd_sc_hd__nor2_2
XFILLER_71_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_5_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7225_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_24_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _5174_/B _5030_/B vssd1 vssd1 vccd1 vccd1 _5032_/A sky130_fd_sc_hd__xor2_2
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7292__85 vssd1 vssd1 vccd1 vccd1 _7292__85/HI _7400_/A sky130_fd_sc_hd__conb_1
X_6981_ _6981_/A _6983_/B vssd1 vssd1 vccd1 vccd1 _6981_/Y sky130_fd_sc_hd__nand2_1
XFILLER_93_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5932_ _5932_/A _5932_/B vssd1 vssd1 vccd1 vccd1 _5935_/A sky130_fd_sc_hd__and2_1
XFILLER_80_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5863_ _5863_/A _5867_/A _5863_/C vssd1 vssd1 vccd1 vccd1 _5864_/B sky130_fd_sc_hd__and3_1
X_4814_ _4814_/A _4814_/B vssd1 vssd1 vccd1 vccd1 _4830_/A sky130_fd_sc_hd__xnor2_1
X_5794_ _6240_/A _6174_/A vssd1 vssd1 vccd1 vccd1 _5795_/B sky130_fd_sc_hd__or2_1
X_4745_ _5749_/A _4745_/B vssd1 vssd1 vccd1 vccd1 _4746_/B sky130_fd_sc_hd__and2_1
X_4676_ _4676_/A _4741_/B vssd1 vssd1 vccd1 vccd1 _4676_/Y sky130_fd_sc_hd__nand2_1
X_7395_ _7395_/A _3689_/Y vssd1 vssd1 vccd1 vccd1 io_out[37] sky130_fd_sc_hd__ebufn_8
X_3627_ _3629_/A vssd1 vssd1 vccd1 vccd1 _3627_/Y sky130_fd_sc_hd__inv_2
X_6415_ _6607_/B _6415_/B vssd1 vssd1 vccd1 vccd1 _6711_/A sky130_fd_sc_hd__and2b_1
X_6346_ _6369_/B _6346_/B _6346_/C vssd1 vssd1 vccd1 vccd1 _6347_/B sky130_fd_sc_hd__nor3_1
XFILLER_88_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6277_ _7006_/A _6132_/Y _6043_/Y vssd1 vssd1 vccd1 vccd1 _6325_/B sky130_fd_sc_hd__a21oi_2
X_5228_ _6045_/B _5228_/B vssd1 vssd1 vccd1 vccd1 _5229_/C sky130_fd_sc_hd__or2_1
X_5159_ _5606_/B vssd1 vssd1 vccd1 vccd1 _6240_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4530_ _4857_/B vssd1 vssd1 vccd1 vccd1 _7078_/A sky130_fd_sc_hd__buf_2
X_4461_ _4470_/B _4469_/C _4469_/B _6410_/A vssd1 vssd1 vccd1 vccd1 _4564_/A sky130_fd_sc_hd__and4b_1
XFILLER_7_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6200_ _6021_/X _6796_/A _6199_/Y vssd1 vssd1 vccd1 vccd1 _6204_/A sky130_fd_sc_hd__a21o_1
X_7180_ _7183_/CLK _7180_/D vssd1 vssd1 vccd1 vccd1 _7180_/Q sky130_fd_sc_hd__dfxtp_1
X_4392_ _7208_/Q _4392_/B vssd1 vssd1 vccd1 vccd1 _4393_/B sky130_fd_sc_hd__or2_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6131_ _6198_/A _6198_/B vssd1 vssd1 vccd1 vccd1 _6217_/A sky130_fd_sc_hd__xnor2_2
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _6063_/A _6063_/B _6063_/C vssd1 vssd1 vccd1 vccd1 _6064_/A sky130_fd_sc_hd__o21a_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5013_ _6140_/A _6136_/A vssd1 vssd1 vccd1 vccd1 _5014_/B sky130_fd_sc_hd__nand2_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6964_ _6977_/A vssd1 vssd1 vccd1 vccd1 _6964_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5915_ _5915_/A _5915_/B vssd1 vssd1 vccd1 vccd1 _5950_/A sky130_fd_sc_hd__or2_1
X_6895_ hold15/X _6892_/X _6894_/X hold51/A vssd1 vssd1 vccd1 vccd1 _6895_/X sky130_fd_sc_hd__a22o_1
XFILLER_42_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5846_ _5865_/A _5865_/B _5845_/X vssd1 vssd1 vccd1 vccd1 _6092_/B sky130_fd_sc_hd__a21oi_2
XFILLER_21_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5777_ _5821_/A _5821_/B vssd1 vssd1 vccd1 vccd1 _5777_/X sky130_fd_sc_hd__and2_1
X_4728_ hold71/A _4728_/B _4728_/C vssd1 vssd1 vccd1 vccd1 _4802_/A sky130_fd_sc_hd__and3_1
X_4659_ _4659_/A _4659_/B vssd1 vssd1 vccd1 vccd1 _4660_/B sky130_fd_sc_hd__nor2_1
XFILLER_101_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7378_ _7378_/A _3668_/Y vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__ebufn_8
XFILLER_88_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6329_ _6329_/A _6329_/B vssd1 vssd1 vccd1 vccd1 _6330_/B sky130_fd_sc_hd__nand2_1
XFILLER_49_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7262__55 vssd1 vssd1 vccd1 vccd1 _7262__55/HI _7361_/A sky130_fd_sc_hd__conb_1
XFILLER_35_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3961_ _3960_/A _4157_/A _4154_/A _3960_/D vssd1 vssd1 vccd1 vccd1 _3962_/B sky130_fd_sc_hd__a22o_1
XFILLER_90_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5700_ _5700_/A _5700_/B vssd1 vssd1 vccd1 vccd1 _5716_/B sky130_fd_sc_hd__xnor2_4
XFILLER_50_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6680_ _6687_/B _6926_/A _6688_/A vssd1 vssd1 vccd1 vccd1 _6681_/A sky130_fd_sc_hd__and3_1
X_3892_ _4951_/A _4951_/B vssd1 vssd1 vccd1 vccd1 _3933_/A sky130_fd_sc_hd__xnor2_1
X_5631_ _5869_/B _5869_/A vssd1 vssd1 vccd1 vccd1 _5631_/X sky130_fd_sc_hd__or2b_1
X_5562_ _5563_/A _5563_/B vssd1 vssd1 vccd1 vccd1 _5564_/A sky130_fd_sc_hd__or2_1
X_4513_ _4514_/A _4514_/B vssd1 vssd1 vccd1 vccd1 _4604_/B sky130_fd_sc_hd__xor2_2
Xhold103 _7196_/Q vssd1 vssd1 vccd1 vccd1 _3825_/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold125 _7033_/A vssd1 vssd1 vccd1 vccd1 hold125/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold114 hold27/X vssd1 vssd1 vccd1 vccd1 hold114/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_5493_ _5493_/A _5538_/B vssd1 vssd1 vccd1 vccd1 _5496_/A sky130_fd_sc_hd__xor2_1
X_4444_ _4444_/A _4444_/B vssd1 vssd1 vccd1 vccd1 _4523_/A sky130_fd_sc_hd__xnor2_1
X_7163_ _7172_/CLK _7163_/D vssd1 vssd1 vccd1 vccd1 _7163_/Q sky130_fd_sc_hd__dfxtp_2
X_4375_ _5719_/A _4375_/B vssd1 vssd1 vccd1 vccd1 _4375_/Y sky130_fd_sc_hd__nor2_1
X_7094_ hold84/X _7088_/X _7093_/Y _7086_/X vssd1 vssd1 vccd1 vccd1 hold86/A sky130_fd_sc_hd__o211a_1
X_6114_ _6796_/A _6114_/B vssd1 vssd1 vccd1 vccd1 _6115_/B sky130_fd_sc_hd__xnor2_2
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6045_ _7001_/A _6045_/B vssd1 vssd1 vccd1 vccd1 _6046_/B sky130_fd_sc_hd__nor2_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6947_ _6947_/A _6956_/B vssd1 vssd1 vccd1 vccd1 _6947_/Y sky130_fd_sc_hd__nand2_1
XFILLER_54_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6878_ _6877_/A _6877_/B _6877_/C vssd1 vssd1 vccd1 vccd1 _6878_/Y sky130_fd_sc_hd__a21oi_1
X_5829_ _7016_/A _5829_/B vssd1 vssd1 vccd1 vccd1 _5829_/X sky130_fd_sc_hd__and2_1
XFILLER_89_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4160_ _4038_/A _4064_/A _4065_/B _4065_/A vssd1 vssd1 vccd1 vccd1 _4162_/B sky130_fd_sc_hd__a22oi_2
XFILLER_95_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4091_ _4097_/B vssd1 vssd1 vccd1 vccd1 _6613_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_82_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6801_ _6983_/A _6825_/B vssd1 vssd1 vccd1 vccd1 _6829_/A sky130_fd_sc_hd__xnor2_1
XFILLER_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4993_ _4993_/A _4993_/B vssd1 vssd1 vccd1 vccd1 _4994_/B sky130_fd_sc_hd__nor2_1
X_3944_ _7214_/Q _3944_/B vssd1 vssd1 vccd1 vccd1 _4189_/A sky130_fd_sc_hd__xnor2_4
X_6732_ _6732_/A _6767_/B vssd1 vssd1 vccd1 vccd1 _6763_/A sky130_fd_sc_hd__nand2_2
X_3875_ _7198_/Q vssd1 vssd1 vccd1 vccd1 _4957_/A sky130_fd_sc_hd__clkbuf_2
X_6663_ _6687_/B _6676_/A _6677_/A vssd1 vssd1 vccd1 vccd1 _6664_/B sky130_fd_sc_hd__o21ai_1
X_5614_ _5614_/A _5614_/B vssd1 vssd1 vccd1 vccd1 _5634_/B sky130_fd_sc_hd__xor2_2
X_6594_ _6593_/B _6594_/B vssd1 vssd1 vccd1 vccd1 _6594_/X sky130_fd_sc_hd__and2b_1
X_5545_ _5508_/A _5507_/B _5507_/A vssd1 vssd1 vccd1 vccd1 _5553_/A sky130_fd_sc_hd__a21bo_1
X_5476_ _5476_/A _5476_/B vssd1 vssd1 vccd1 vccd1 _5526_/A sky130_fd_sc_hd__nor2_1
X_4427_ _4543_/A _4543_/B vssd1 vssd1 vccd1 vccd1 _4641_/A sky130_fd_sc_hd__and2_2
X_7215_ _7222_/CLK _7215_/D vssd1 vssd1 vccd1 vccd1 _7215_/Q sky130_fd_sc_hd__dfxtp_1
X_7146_ _7226_/CLK _7146_/D vssd1 vssd1 vccd1 vccd1 _7385_/A sky130_fd_sc_hd__dfxtp_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4358_ hold53/X vssd1 vssd1 vccd1 vccd1 _7070_/A sky130_fd_sc_hd__inv_2
X_7077_ _5478_/A _7075_/X _7076_/X _7073_/X vssd1 vssd1 vccd1 vccd1 _7207_/D sky130_fd_sc_hd__o211a_1
XFILLER_58_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4289_ _4289_/A _4289_/B vssd1 vssd1 vccd1 vccd1 _4291_/B sky130_fd_sc_hd__xor2_1
XFILLER_86_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6028_ _7191_/Q _7025_/A vssd1 vssd1 vccd1 vccd1 _6118_/B sky130_fd_sc_hd__xnor2_2
XFILLER_64_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7232__25 vssd1 vssd1 vccd1 vccd1 _7232__25/HI _7331_/A sky130_fd_sc_hd__conb_1
XFILLER_33_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3660_ _3660_/A vssd1 vssd1 vccd1 vccd1 _3660_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5330_ _5330_/A vssd1 vssd1 vccd1 vccd1 _5330_/Y sky130_fd_sc_hd__inv_2
X_5261_ hold74/X vssd1 vssd1 vccd1 vccd1 _6261_/A sky130_fd_sc_hd__buf_2
X_4212_ _7089_/A _4856_/A hold71/A vssd1 vssd1 vccd1 vccd1 _4408_/B sky130_fd_sc_hd__o21ai_1
X_7000_ _6975_/A _6993_/X _6999_/Y _6995_/X vssd1 vssd1 vccd1 vccd1 _7178_/D sky130_fd_sc_hd__o211a_1
X_5192_ _7173_/Q vssd1 vssd1 vccd1 vccd1 _6546_/A sky130_fd_sc_hd__clkbuf_1
X_4143_ _5783_/B _5168_/A _6617_/A _6063_/A vssd1 vssd1 vccd1 vccd1 _4143_/X sky130_fd_sc_hd__a31o_1
XFILLER_95_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4074_ _6483_/B vssd1 vssd1 vccd1 vccd1 _4721_/A sky130_fd_sc_hd__inv_2
XFILLER_55_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7311__104 vssd1 vssd1 vccd1 vccd1 _7311__104/HI _7419_/A sky130_fd_sc_hd__conb_1
XFILLER_24_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4976_ _5118_/A _5118_/B vssd1 vssd1 vccd1 vccd1 _4978_/C sky130_fd_sc_hd__xnor2_1
XFILLER_11_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6715_ _6758_/B _6715_/B vssd1 vssd1 vccd1 vccd1 _6716_/B sky130_fd_sc_hd__and2b_1
X_3927_ _3928_/B _3927_/B vssd1 vssd1 vccd1 vccd1 _4008_/B sky130_fd_sc_hd__xnor2_1
X_3858_ _4252_/A _3848_/Y _3920_/A _3857_/Y vssd1 vssd1 vccd1 vccd1 _4950_/B sky130_fd_sc_hd__o22ai_4
X_6646_ _6649_/A _6649_/B _6645_/X vssd1 vssd1 vccd1 vccd1 _6647_/B sky130_fd_sc_hd__a21oi_2
X_3789_ hold98/A _4356_/B vssd1 vssd1 vccd1 vccd1 _5056_/B sky130_fd_sc_hd__or2_1
X_6577_ _6577_/A _6600_/B vssd1 vssd1 vccd1 vccd1 _6603_/A sky130_fd_sc_hd__nor2_1
X_5528_ _5528_/A _5467_/B vssd1 vssd1 vccd1 vccd1 _5529_/B sky130_fd_sc_hd__or2b_1
XFILLER_3_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5459_ _5360_/A _5360_/B _5322_/A vssd1 vssd1 vccd1 vccd1 _5521_/B sky130_fd_sc_hd__a21oi_1
X_7298__91 vssd1 vssd1 vccd1 vccd1 _7298__91/HI _7406_/A sky130_fd_sc_hd__conb_1
XFILLER_101_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7129_ _7151_/CLK _7129_/D vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__dfxtp_1
XFILLER_19_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4830_ _4830_/A _4830_/B vssd1 vssd1 vccd1 vccd1 _4927_/A sky130_fd_sc_hd__nor2_1
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4761_ _4761_/A _4761_/B vssd1 vssd1 vccd1 vccd1 _4772_/A sky130_fd_sc_hd__xor2_2
X_3712_ _3715_/A vssd1 vssd1 vccd1 vccd1 _3712_/Y sky130_fd_sc_hd__inv_2
X_4692_ _4692_/A _4692_/B vssd1 vssd1 vccd1 vccd1 _4707_/A sky130_fd_sc_hd__xnor2_2
X_6500_ _6487_/X _6497_/Y _6493_/X _6505_/A vssd1 vssd1 vccd1 vccd1 _6506_/B sky130_fd_sc_hd__o211ai_1
X_6431_ _6484_/A _6483_/A _6485_/B vssd1 vssd1 vccd1 vccd1 _6432_/C sky130_fd_sc_hd__nand3_1
X_3643_ _3647_/A vssd1 vssd1 vccd1 vccd1 _3643_/Y sky130_fd_sc_hd__inv_2
X_6362_ _6335_/A _6362_/B vssd1 vssd1 vccd1 vccd1 _6365_/B sky130_fd_sc_hd__and2b_1
X_5313_ _6270_/A _5483_/C vssd1 vssd1 vccd1 vccd1 _5314_/B sky130_fd_sc_hd__xor2_2
XFILLER_88_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6293_ _6294_/B _6293_/B vssd1 vssd1 vccd1 vccd1 _6295_/A sky130_fd_sc_hd__and2b_1
XFILLER_88_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5244_ _5096_/A _5096_/B _5243_/X vssd1 vssd1 vccd1 vccd1 _5368_/B sky130_fd_sc_hd__a21bo_1
X_5175_ _5029_/A _5029_/B _5174_/X vssd1 vssd1 vccd1 vccd1 _5176_/B sky130_fd_sc_hd__a21oi_4
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_4126_ _7182_/Q vssd1 vssd1 vccd1 vccd1 _4374_/A sky130_fd_sc_hd__clkbuf_1
X_4057_ _6016_/A vssd1 vssd1 vccd1 vccd1 _6449_/A sky130_fd_sc_hd__inv_2
XFILLER_56_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4959_ _5277_/B _4959_/B vssd1 vssd1 vccd1 vccd1 _5286_/A sky130_fd_sc_hd__or2_1
XFILLER_61_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6629_ _6973_/A _6655_/B vssd1 vssd1 vccd1 vccd1 _6656_/A sky130_fd_sc_hd__nor2_1
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6980_ _6794_/A _6977_/X _6978_/Y _6979_/X vssd1 vssd1 vccd1 vccd1 _7171_/D sky130_fd_sc_hd__o211a_1
XFILLER_93_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5931_ _5931_/A vssd1 vssd1 vccd1 vccd1 _5932_/B sky130_fd_sc_hd__clkinv_2
XFILLER_18_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5862_ _5862_/A _5862_/B vssd1 vssd1 vccd1 vccd1 _6097_/A sky130_fd_sc_hd__xnor2_2
X_4813_ _4865_/A _4813_/B vssd1 vssd1 vccd1 vccd1 _4928_/A sky130_fd_sc_hd__xnor2_1
XFILLER_33_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5793_ _6076_/A _5793_/B vssd1 vssd1 vccd1 vccd1 _5798_/A sky130_fd_sc_hd__or2_1
X_4744_ _6409_/A _4744_/B vssd1 vssd1 vccd1 vccd1 _4790_/A sky130_fd_sc_hd__nand2_2
X_4675_ _6137_/B _5749_/A _5812_/A vssd1 vssd1 vccd1 vccd1 _4742_/B sky130_fd_sc_hd__or3_1
X_7394_ _7394_/A _3688_/Y vssd1 vssd1 vccd1 vccd1 io_out[36] sky130_fd_sc_hd__ebufn_8
X_6414_ _6413_/A _4092_/Y _6584_/A vssd1 vssd1 vccd1 vccd1 _6415_/B sky130_fd_sc_hd__a21o_1
X_3626_ _3629_/A vssd1 vssd1 vccd1 vccd1 _3626_/Y sky130_fd_sc_hd__inv_2
X_6345_ _6346_/B _6346_/C _6369_/B vssd1 vssd1 vccd1 vccd1 _6383_/A sky130_fd_sc_hd__o21a_1
X_6276_ _6324_/A _6276_/B vssd1 vssd1 vccd1 vccd1 _6325_/A sky130_fd_sc_hd__xnor2_2
X_7268__61 vssd1 vssd1 vccd1 vccd1 _7268__61/HI _7367_/A sky130_fd_sc_hd__conb_1
X_5227_ _5406_/A _6132_/A vssd1 vssd1 vccd1 vccd1 _5229_/B sky130_fd_sc_hd__nand2_1
XFILLER_88_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5158_ _4994_/A _4994_/B _4993_/A vssd1 vssd1 vccd1 vccd1 _5325_/A sky130_fd_sc_hd__a21o_1
XFILLER_29_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7317__110 vssd1 vssd1 vccd1 vccd1 _7317__110/HI _7425_/A sky130_fd_sc_hd__conb_1
XFILLER_56_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4109_ _7165_/Q _5021_/A _7166_/Q vssd1 vssd1 vccd1 vccd1 _4138_/B sky130_fd_sc_hd__a21oi_4
XFILLER_17_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5089_ _4384_/A _4384_/B _4383_/A vssd1 vssd1 vccd1 vccd1 _5091_/B sky130_fd_sc_hd__a21oi_2
XFILLER_71_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4460_ _4460_/A vssd1 vssd1 vccd1 vccd1 _6410_/A sky130_fd_sc_hd__buf_2
XFILLER_7_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4391_ _4391_/A _4391_/B vssd1 vssd1 vccd1 vccd1 _4522_/A sky130_fd_sc_hd__xnor2_4
X_6130_ _6033_/A _6128_/X _6124_/A _6129_/Y vssd1 vssd1 vccd1 vccd1 _6198_/B sky130_fd_sc_hd__o31a_1
XFILLER_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _6174_/A _6061_/B vssd1 vssd1 vccd1 vccd1 _6063_/C sky130_fd_sc_hd__xor2_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _5762_/A vssd1 vssd1 vccd1 vccd1 _6136_/A sky130_fd_sc_hd__clkinv_2
XFILLER_66_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6963_ _4429_/A _6949_/X _6962_/X _6952_/X vssd1 vssd1 vccd1 vccd1 _7165_/D sky130_fd_sc_hd__o211a_1
X_5914_ _5914_/A _5914_/B vssd1 vssd1 vccd1 vccd1 _5915_/B sky130_fd_sc_hd__and2_1
X_6894_ _6894_/A vssd1 vssd1 vccd1 vccd1 _6894_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5845_ _5844_/B _5845_/B vssd1 vssd1 vccd1 vccd1 _5845_/X sky130_fd_sc_hd__and2b_1
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5776_ _5761_/Y _5774_/B _5775_/Y vssd1 vssd1 vccd1 vccd1 _5821_/B sky130_fd_sc_hd__o21a_1
X_4727_ _4799_/A _4857_/B _4412_/A vssd1 vssd1 vccd1 vccd1 _4728_/C sky130_fd_sc_hd__o21ai_1
XFILLER_21_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4658_ _4658_/A _4658_/B vssd1 vssd1 vccd1 vccd1 _4733_/B sky130_fd_sc_hd__or2_1
X_3609_ input1/X vssd1 vssd1 vccd1 vccd1 _3734_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_89_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4589_ _6625_/A vssd1 vssd1 vccd1 vccd1 _6620_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7377_ _7377_/A _3666_/Y vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__ebufn_8
XFILLER_88_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6328_ _6329_/A _6329_/B vssd1 vssd1 vccd1 vccd1 _6330_/A sky130_fd_sc_hd__or2_1
XFILLER_88_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6259_ _6257_/X _6258_/Y _6261_/A vssd1 vssd1 vccd1 vccd1 _6259_/X sky130_fd_sc_hd__a21o_1
XFILLER_76_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3960_ _3960_/A _4157_/A _4154_/A _3960_/D vssd1 vssd1 vccd1 vccd1 _4157_/B sky130_fd_sc_hd__nand4_2
XFILLER_63_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3891_ _4981_/A _3891_/B vssd1 vssd1 vccd1 vccd1 _4951_/B sky130_fd_sc_hd__xnor2_1
X_5630_ _5630_/A _5812_/B vssd1 vssd1 vccd1 vccd1 _5869_/A sky130_fd_sc_hd__xor2_2
X_5561_ _5520_/A _5520_/B _5560_/X vssd1 vssd1 vccd1 vccd1 _5563_/B sky130_fd_sc_hd__o21a_1
X_4512_ _4499_/Y _4607_/B _4511_/Y vssd1 vssd1 vccd1 vccd1 _4514_/B sky130_fd_sc_hd__a21o_1
X_5492_ _5546_/A _5492_/B vssd1 vssd1 vccd1 vccd1 _5538_/B sky130_fd_sc_hd__xnor2_1
Xhold104 _3770_/A vssd1 vssd1 vccd1 vccd1 _7028_/A sky130_fd_sc_hd__clkbuf_2
Xhold115 hold40/X vssd1 vssd1 vccd1 vccd1 _3746_/B sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold126 _6104_/X vssd1 vssd1 vccd1 vccd1 hold126/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4443_ _4443_/A _4443_/B vssd1 vssd1 vccd1 vccd1 _4444_/B sky130_fd_sc_hd__and2_2
X_7162_ _7172_/CLK _7162_/D vssd1 vssd1 vccd1 vccd1 _7162_/Q sky130_fd_sc_hd__dfxtp_2
X_4374_ _4374_/A vssd1 vssd1 vccd1 vccd1 _5719_/A sky130_fd_sc_hd__clkbuf_4
X_7093_ _7093_/A _7093_/B vssd1 vssd1 vccd1 vccd1 _7093_/Y sky130_fd_sc_hd__nand2_1
X_6113_ _6470_/A _6938_/A _6021_/X vssd1 vssd1 vccd1 vccd1 _6114_/B sky130_fd_sc_hd__a21oi_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7238__31 vssd1 vssd1 vccd1 vccd1 _7238__31/HI _7337_/A sky130_fd_sc_hd__conb_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6044_ _6136_/A _6043_/Y _7001_/A vssd1 vssd1 vccd1 vccd1 _6046_/A sky130_fd_sc_hd__mux2_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6946_ input8/X _6935_/X _6945_/Y _6939_/X vssd1 vssd1 vccd1 vccd1 _7159_/D sky130_fd_sc_hd__o211a_1
XFILLER_54_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6877_ _6877_/A _6877_/B _6877_/C vssd1 vssd1 vccd1 vccd1 _6877_/X sky130_fd_sc_hd__and3_1
X_5828_ _7016_/A _5829_/B vssd1 vssd1 vccd1 vccd1 _5872_/B sky130_fd_sc_hd__xor2_2
XFILLER_22_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5759_ _5759_/A _5759_/B vssd1 vssd1 vccd1 vccd1 _5821_/A sky130_fd_sc_hd__xnor2_2
X_7429_ _7429_/A _3727_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[33] sky130_fd_sc_hd__ebufn_8
XFILLER_78_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4090_ _7165_/Q _7164_/Q vssd1 vssd1 vccd1 vccd1 _4097_/B sky130_fd_sc_hd__xor2_4
XFILLER_36_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6800_ _6824_/A _6824_/B vssd1 vssd1 vccd1 vccd1 _6825_/B sky130_fd_sc_hd__xnor2_1
XFILLER_36_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4992_ _4992_/A _4992_/B _4992_/C vssd1 vssd1 vccd1 vccd1 _4993_/B sky130_fd_sc_hd__and3_1
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3943_ _4026_/A _3943_/B vssd1 vssd1 vccd1 vccd1 _3963_/A sky130_fd_sc_hd__xor2_1
X_6731_ _6730_/A _6730_/B _6730_/C vssd1 vssd1 vccd1 vccd1 _6767_/B sky130_fd_sc_hd__a21o_1
XFILLER_16_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3874_ _4003_/A vssd1 vssd1 vccd1 vccd1 _3879_/B sky130_fd_sc_hd__buf_2
X_6662_ _6662_/A _6662_/B vssd1 vssd1 vccd1 vccd1 _6677_/A sky130_fd_sc_hd__nand2_1
X_5613_ _5801_/B _5613_/B vssd1 vssd1 vccd1 vccd1 _5614_/B sky130_fd_sc_hd__xor2_2
X_6593_ _6594_/B _6593_/B vssd1 vssd1 vccd1 vccd1 _6620_/B sky130_fd_sc_hd__xnor2_2
X_5544_ _5584_/A _5584_/B vssd1 vssd1 vccd1 vccd1 _5554_/A sky130_fd_sc_hd__xnor2_1
X_5475_ _5475_/A _5475_/B vssd1 vssd1 vccd1 vccd1 _5531_/A sky130_fd_sc_hd__nand2_1
X_4426_ _4426_/A _7217_/Q vssd1 vssd1 vccd1 vccd1 _4543_/B sky130_fd_sc_hd__xnor2_1
X_7214_ _7222_/CLK hold86/X vssd1 vssd1 vccd1 vccd1 _7214_/Q sky130_fd_sc_hd__dfxtp_2
X_7145_ _7151_/CLK hold33/X vssd1 vssd1 vccd1 vccd1 _7384_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_86_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4357_ hold85/A hold59/A vssd1 vssd1 vccd1 vccd1 _5062_/C sky130_fd_sc_hd__xor2_1
XFILLER_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7076_ hold82/X _7091_/B vssd1 vssd1 vccd1 vccd1 _7076_/X sky130_fd_sc_hd__or2_1
XFILLER_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4288_ _6039_/B _6045_/B _5827_/A vssd1 vssd1 vccd1 vccd1 _4289_/B sky130_fd_sc_hd__mux2_1
X_6027_ _6027_/A vssd1 vssd1 vccd1 vccd1 _7025_/A sky130_fd_sc_hd__buf_2
XFILLER_73_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6929_ _6929_/A _6933_/B vssd1 vssd1 vccd1 vccd1 _6929_/Y sky130_fd_sc_hd__nand2_1
XFILLER_80_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_49_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5260_ _3750_/X hold19/X _3752_/X _5259_/X vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__o211a_1
X_4211_ _7217_/Q vssd1 vssd1 vccd1 vccd1 _4856_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5191_ _5198_/B vssd1 vssd1 vccd1 vccd1 _6564_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_95_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4142_ _7167_/Q _5006_/B vssd1 vssd1 vccd1 vccd1 _6063_/A sky130_fd_sc_hd__and2_1
X_4073_ _6485_/B vssd1 vssd1 vccd1 vccd1 _6483_/B sky130_fd_sc_hd__buf_2
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4975_ _4975_/A _5148_/B vssd1 vssd1 vccd1 vccd1 _5118_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3926_ _3844_/X _4506_/C _4009_/B vssd1 vssd1 vccd1 vccd1 _3927_/B sky130_fd_sc_hd__a21boi_1
X_6714_ _6715_/B _6758_/B vssd1 vssd1 vccd1 vccd1 _6793_/A sky130_fd_sc_hd__and2b_1
XFILLER_32_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3857_ _7016_/A _3838_/Y _5267_/A _5765_/A vssd1 vssd1 vccd1 vccd1 _3857_/Y sky130_fd_sc_hd__a211oi_2
X_6645_ _6644_/B _6645_/B vssd1 vssd1 vccd1 vccd1 _6645_/X sky130_fd_sc_hd__and2b_1
X_3788_ hold59/X vssd1 vssd1 vccd1 vccd1 hold58/A sky130_fd_sc_hd__clkbuf_2
X_6576_ _6576_/A _6576_/B vssd1 vssd1 vccd1 vccd1 _6600_/B sky130_fd_sc_hd__xnor2_1
X_5527_ _5527_/A _5466_/A vssd1 vssd1 vccd1 vccd1 _5529_/A sky130_fd_sc_hd__or2b_1
X_5458_ _5458_/A _5458_/B vssd1 vssd1 vccd1 vccd1 _5521_/A sky130_fd_sc_hd__xnor2_1
XFILLER_99_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4409_ _4409_/A _4409_/B vssd1 vssd1 vccd1 vccd1 _4538_/A sky130_fd_sc_hd__xnor2_2
X_5389_ _7091_/A _6945_/A vssd1 vssd1 vccd1 vccd1 _5397_/B sky130_fd_sc_hd__nand2_1
XFILLER_59_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7128_ _7151_/CLK hold29/X vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__dfxtp_1
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7059_ hold70/X _7059_/B vssd1 vssd1 vccd1 vccd1 _7059_/X sky130_fd_sc_hd__or2_1
XFILLER_59_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4760_ _4760_/A _4760_/B vssd1 vssd1 vccd1 vccd1 _4775_/A sky130_fd_sc_hd__xnor2_2
XFILLER_81_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4691_ _4691_/A _4734_/A vssd1 vssd1 vccd1 vccd1 _4758_/A sky130_fd_sc_hd__xor2_1
X_3711_ _3715_/A vssd1 vssd1 vccd1 vccd1 _3711_/Y sky130_fd_sc_hd__inv_2
X_3642_ _3648_/A vssd1 vssd1 vccd1 vccd1 _3647_/A sky130_fd_sc_hd__buf_12
X_6430_ _6494_/A _6485_/B _7157_/Q vssd1 vssd1 vccd1 vccd1 _6432_/B sky130_fd_sc_hd__a21o_1
X_6361_ _6261_/X _6359_/X _6360_/X _6196_/X vssd1 vssd1 vccd1 vccd1 _7133_/D sky130_fd_sc_hd__o211a_1
X_5312_ _5406_/A _6966_/A vssd1 vssd1 vccd1 vccd1 _5483_/C sky130_fd_sc_hd__nand2_2
X_6292_ _6346_/B _6292_/B vssd1 vssd1 vccd1 vccd1 _6293_/B sky130_fd_sc_hd__or2_1
X_5243_ _5243_/A _5041_/B vssd1 vssd1 vccd1 vccd1 _5243_/X sky130_fd_sc_hd__or2b_1
X_5174_ _5030_/B _5174_/B vssd1 vssd1 vccd1 vccd1 _5174_/X sky130_fd_sc_hd__and2b_1
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4125_ _7182_/Q _5011_/A vssd1 vssd1 vccd1 vccd1 _4286_/A sky130_fd_sc_hd__nand2_1
XFILLER_56_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4056_ _4795_/A vssd1 vssd1 vccd1 vccd1 _4794_/A sky130_fd_sc_hd__buf_2
XFILLER_45_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4958_ _5121_/A _4957_/C _5276_/A vssd1 vssd1 vccd1 vccd1 _4959_/B sky130_fd_sc_hd__a21oi_1
X_4889_ _4889_/A _4889_/B vssd1 vssd1 vccd1 vccd1 _4890_/B sky130_fd_sc_hd__and2_1
X_3909_ _3965_/A _3909_/B vssd1 vssd1 vccd1 vccd1 _3918_/A sky130_fd_sc_hd__xnor2_1
X_6628_ _6628_/A _6628_/B vssd1 vssd1 vccd1 vccd1 _6655_/B sky130_fd_sc_hd__xnor2_1
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6559_ _6559_/A _6410_/A vssd1 vssd1 vccd1 vccd1 _6559_/X sky130_fd_sc_hd__or2b_1
XFILLER_3_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5930_ _5930_/A _5930_/B vssd1 vssd1 vccd1 vccd1 _5935_/B sky130_fd_sc_hd__xor2_1
XFILLER_18_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5861_ _5861_/A _5861_/B vssd1 vssd1 vccd1 vccd1 _5862_/B sky130_fd_sc_hd__xor2_2
X_4812_ _4812_/A _4812_/B vssd1 vssd1 vccd1 vccd1 _4833_/B sky130_fd_sc_hd__xor2_1
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5792_ _5792_/A _5792_/B vssd1 vssd1 vccd1 vccd1 _5793_/B sky130_fd_sc_hd__nor2_1
XFILLER_21_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4743_ _5597_/B vssd1 vssd1 vccd1 vccd1 _6409_/A sky130_fd_sc_hd__clkbuf_2
X_4674_ _4674_/A vssd1 vssd1 vccd1 vccd1 _5749_/A sky130_fd_sc_hd__clkbuf_2
X_6413_ _6413_/A _6413_/B vssd1 vssd1 vccd1 vccd1 _6584_/A sky130_fd_sc_hd__nor2_1
X_3625_ _3629_/A vssd1 vssd1 vccd1 vccd1 _3625_/Y sky130_fd_sc_hd__inv_2
X_7393_ _7393_/A _3687_/Y vssd1 vssd1 vccd1 vccd1 io_out[35] sky130_fd_sc_hd__ebufn_8
X_6344_ _6344_/A _6380_/B vssd1 vssd1 vccd1 vccd1 _6348_/A sky130_fd_sc_hd__xor2_1
XFILLER_88_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6275_ _6327_/A _6324_/C vssd1 vssd1 vccd1 vccd1 _6276_/B sky130_fd_sc_hd__and2_1
XFILLER_88_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5226_ _6139_/A _5226_/B vssd1 vssd1 vccd1 vccd1 _6132_/A sky130_fd_sc_hd__nor2_2
XFILLER_56_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5157_ _5032_/A _5032_/B _5156_/X vssd1 vssd1 vccd1 vccd1 _5181_/A sky130_fd_sc_hd__o21ai_4
X_4108_ _4279_/A _5021_/A vssd1 vssd1 vccd1 vccd1 _4110_/A sky130_fd_sc_hd__nor2_1
X_7283__76 vssd1 vssd1 vccd1 vccd1 _7283__76/HI _7382_/A sky130_fd_sc_hd__conb_1
XFILLER_29_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5088_ _5088_/A _5088_/B vssd1 vssd1 vccd1 vccd1 _5091_/A sky130_fd_sc_hd__xnor2_2
X_4039_ _4039_/A _4039_/B vssd1 vssd1 vccd1 vccd1 _4039_/X sky130_fd_sc_hd__and2_1
XFILLER_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4390_ _5101_/B _4390_/B vssd1 vssd1 vccd1 vccd1 _4391_/B sky130_fd_sc_hd__xnor2_4
XFILLER_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ _5744_/A _5744_/B _5747_/B vssd1 vssd1 vccd1 vccd1 _6075_/A sky130_fd_sc_hd__a21bo_1
XFILLER_85_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _5011_/A vssd1 vssd1 vccd1 vccd1 _5762_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_66_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6962_ _6962_/A _6975_/B vssd1 vssd1 vccd1 vccd1 _6962_/X sky130_fd_sc_hd__or2_1
X_5913_ _5913_/A _5913_/B vssd1 vssd1 vccd1 vccd1 _5944_/B sky130_fd_sc_hd__xnor2_2
X_6893_ _6893_/A _6893_/B vssd1 vssd1 vccd1 vccd1 _6894_/A sky130_fd_sc_hd__nor2_1
XFILLER_34_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5844_ _5845_/B _5844_/B vssd1 vssd1 vccd1 vccd1 _5865_/B sky130_fd_sc_hd__xnor2_1
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5775_ _5840_/A _5840_/B vssd1 vssd1 vccd1 vccd1 _5775_/Y sky130_fd_sc_hd__nand2_1
X_4726_ _4799_/B _4726_/B vssd1 vssd1 vccd1 vccd1 _4728_/B sky130_fd_sc_hd__or2_1
X_4657_ _4657_/A _4666_/B vssd1 vssd1 vccd1 vccd1 _4658_/B sky130_fd_sc_hd__and2_1
X_7376_ _7376_/A _3665_/Y vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__ebufn_8
X_4588_ _6624_/A vssd1 vssd1 vccd1 vccd1 _6625_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6327_ _6327_/A _6327_/B vssd1 vssd1 vccd1 vccd1 _6329_/B sky130_fd_sc_hd__xnor2_1
X_6258_ _6258_/A _6258_/B vssd1 vssd1 vccd1 vccd1 _6258_/Y sky130_fd_sc_hd__nand2_1
X_5209_ hold58/A _5209_/B vssd1 vssd1 vccd1 vccd1 _5210_/B sky130_fd_sc_hd__or2_1
X_6189_ _6189_/A _6189_/B vssd1 vssd1 vccd1 vccd1 _6189_/X sky130_fd_sc_hd__or2_1
XFILLER_57_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3890_ _4992_/A _3890_/B vssd1 vssd1 vccd1 vccd1 _3891_/B sky130_fd_sc_hd__and2_1
XFILLER_31_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5560_ _5560_/A _5560_/B vssd1 vssd1 vccd1 vccd1 _5560_/X sky130_fd_sc_hd__or2_1
X_4511_ _4511_/A _4511_/B vssd1 vssd1 vccd1 vccd1 _4511_/Y sky130_fd_sc_hd__nor2_1
X_5491_ _5551_/A _5491_/B vssd1 vssd1 vccd1 vccd1 _5492_/B sky130_fd_sc_hd__and2_1
Xhold116 _7041_/A vssd1 vssd1 vccd1 vccd1 hold116/X sky130_fd_sc_hd__clkbuf_1
X_4442_ _4442_/A _4442_/B vssd1 vssd1 vccd1 vccd1 _4443_/B sky130_fd_sc_hd__or2_1
Xhold105 _6120_/B vssd1 vssd1 vccd1 vccd1 _3754_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold127 _7038_/A vssd1 vssd1 vccd1 vccd1 hold127/X sky130_fd_sc_hd__dlygate4sd3_1
X_7161_ _7172_/CLK _7161_/D vssd1 vssd1 vccd1 vccd1 _7161_/Q sky130_fd_sc_hd__dfxtp_2
X_4373_ _4379_/A vssd1 vssd1 vccd1 vccd1 _5229_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_98_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7092_ hold122/X _7088_/X _7091_/X _7086_/X vssd1 vssd1 vccd1 vccd1 hold54/A sky130_fd_sc_hd__o211a_1
X_6112_ _6112_/A vssd1 vssd1 vccd1 vccd1 _6796_/A sky130_fd_sc_hd__clkinv_2
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6043_ _6140_/A _6136_/A vssd1 vssd1 vccd1 vccd1 _6043_/Y sky130_fd_sc_hd__nor2_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7253__46 vssd1 vssd1 vccd1 vccd1 _7253__46/HI _7352_/A sky130_fd_sc_hd__conb_1
XFILLER_26_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6945_ _6945_/A _6956_/B vssd1 vssd1 vccd1 vccd1 _6945_/Y sky130_fd_sc_hd__nand2_1
XFILLER_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_81_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6876_ _6876_/A _6876_/B vssd1 vssd1 vccd1 vccd1 _6877_/C sky130_fd_sc_hd__xnor2_1
X_5827_ _5827_/A _5827_/B vssd1 vssd1 vccd1 vccd1 _5833_/A sky130_fd_sc_hd__xnor2_1
X_5758_ _5758_/A _5838_/B vssd1 vssd1 vccd1 vccd1 _5822_/A sky130_fd_sc_hd__xnor2_1
X_4709_ _4758_/A _4758_/B _4708_/X vssd1 vssd1 vccd1 vccd1 _4711_/B sky130_fd_sc_hd__a21o_1
X_5689_ _5689_/A _6531_/A vssd1 vssd1 vccd1 vccd1 _5715_/A sky130_fd_sc_hd__nand2_2
X_7428_ _7428_/A _3726_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[32] sky130_fd_sc_hd__ebufn_8
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7359_ _7359_/A _3646_/Y vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__ebufn_8
XFILLER_89_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6730_ _6730_/A _6730_/B _6730_/C vssd1 vssd1 vccd1 vccd1 _6732_/A sky130_fd_sc_hd__nand3_1
X_4991_ _4992_/A _4992_/B _4992_/C vssd1 vssd1 vccd1 vccd1 _4993_/A sky130_fd_sc_hd__a21oi_1
XFILLER_23_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3942_ _3942_/A _3978_/B vssd1 vssd1 vccd1 vccd1 _3943_/B sky130_fd_sc_hd__or2_1
XFILLER_51_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6661_ _6662_/A _6662_/B vssd1 vssd1 vccd1 vccd1 _6676_/A sky130_fd_sc_hd__nor2_1
X_3873_ _3873_/A _3873_/B vssd1 vssd1 vccd1 vccd1 _3889_/A sky130_fd_sc_hd__nor2_1
X_5612_ _5801_/A _5636_/A vssd1 vssd1 vccd1 vccd1 _5613_/B sky130_fd_sc_hd__or2_1
X_6592_ _6978_/A _6592_/B vssd1 vssd1 vccd1 vccd1 _6593_/B sky130_fd_sc_hd__xnor2_1
X_5543_ _5543_/A _5543_/B vssd1 vssd1 vccd1 vccd1 _5584_/B sky130_fd_sc_hd__xnor2_1
X_5474_ _3750_/X hold118/X _3752_/X _5473_/X vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__o211a_1
X_4425_ _7220_/Q _6502_/B vssd1 vssd1 vccd1 vccd1 _4543_/A sky130_fd_sc_hd__xnor2_1
X_7213_ _7222_/CLK hold54/X vssd1 vssd1 vccd1 vccd1 _7213_/Q sky130_fd_sc_hd__dfxtp_2
X_4356_ _7066_/A _4356_/B _4359_/B vssd1 vssd1 vccd1 vccd1 _5055_/A sky130_fd_sc_hd__or3_1
X_7144_ _7226_/CLK hold38/X vssd1 vssd1 vccd1 vccd1 _7383_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_98_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7075_ _7101_/A vssd1 vssd1 vccd1 vccd1 _7075_/X sky130_fd_sc_hd__clkbuf_2
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4287_ _7180_/Q vssd1 vssd1 vccd1 vccd1 _5827_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_74_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6026_ _5673_/A _6029_/B _5679_/B _5685_/A vssd1 vssd1 vccd1 vccd1 _6128_/B sky130_fd_sc_hd__a2bb2oi_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6928_ _7052_/A vssd1 vssd1 vccd1 vccd1 _6933_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6859_ _6859_/A _6859_/B vssd1 vssd1 vccd1 vccd1 _6860_/B sky130_fd_sc_hd__or2_1
XFILLER_13_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4210_ _4215_/A _4210_/B vssd1 vssd1 vccd1 vccd1 _4409_/A sky130_fd_sc_hd__nor2_2
X_5190_ _5190_/A _5190_/B vssd1 vssd1 vccd1 vccd1 _5200_/A sky130_fd_sc_hd__nand2_1
XFILLER_95_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4141_ _5783_/B _5006_/B vssd1 vssd1 vccd1 vccd1 _6063_/B sky130_fd_sc_hd__nor2_1
X_4072_ _7155_/Q vssd1 vssd1 vccd1 vccd1 _6485_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_91_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4974_ _4974_/A _4974_/B vssd1 vssd1 vccd1 vccd1 _5148_/B sky130_fd_sc_hd__nand2_1
X_3925_ _4613_/A _5267_/A vssd1 vssd1 vccd1 vccd1 _4009_/B sky130_fd_sc_hd__nand2_1
X_6713_ _6713_/A vssd1 vssd1 vccd1 vccd1 _6758_/B sky130_fd_sc_hd__clkbuf_2
X_6644_ _6645_/B _6644_/B vssd1 vssd1 vccd1 vccd1 _6649_/B sky130_fd_sc_hd__xnor2_1
X_3856_ _4526_/B vssd1 vssd1 vccd1 vccd1 _7016_/A sky130_fd_sc_hd__clkbuf_4
X_6575_ _6575_/A _6575_/B vssd1 vssd1 vccd1 vccd1 _6576_/B sky130_fd_sc_hd__xor2_2
X_3787_ _4353_/A _3787_/B vssd1 vssd1 vccd1 vccd1 _4344_/A sky130_fd_sc_hd__or2_2
X_5526_ _5526_/A _5526_/B vssd1 vssd1 vccd1 vccd1 _5530_/A sky130_fd_sc_hd__xnor2_1
X_5457_ _5457_/A _5518_/A vssd1 vssd1 vccd1 vccd1 _5458_/B sky130_fd_sc_hd__xnor2_1
X_4408_ _4408_/A _4408_/B vssd1 vssd1 vccd1 vccd1 _4409_/B sky130_fd_sc_hd__and2_1
XFILLER_59_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5388_ _5391_/A vssd1 vssd1 vccd1 vccd1 _7096_/A sky130_fd_sc_hd__buf_2
X_4339_ _4339_/A _4339_/B vssd1 vssd1 vccd1 vccd1 _4442_/B sky130_fd_sc_hd__xnor2_1
X_7127_ _7226_/CLK hold76/X vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__dfxtp_1
X_7058_ hold120/X _7045_/X _7057_/X _7048_/X vssd1 vssd1 vccd1 vccd1 _7200_/D sky130_fd_sc_hd__o211a_1
XFILLER_86_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6009_ _6009_/A _6009_/B _6009_/C vssd1 vssd1 vccd1 vccd1 _6011_/B sky130_fd_sc_hd__and3_2
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7289__82 vssd1 vssd1 vccd1 vccd1 _7289__82/HI _7397_/A sky130_fd_sc_hd__conb_1
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3710_ _3710_/A vssd1 vssd1 vccd1 vccd1 _3715_/A sky130_fd_sc_hd__buf_12
X_4690_ _4690_/A _4690_/B vssd1 vssd1 vccd1 vccd1 _4710_/A sky130_fd_sc_hd__xnor2_1
X_3641_ _3641_/A vssd1 vssd1 vccd1 vccd1 _3641_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6360_ _6391_/A hold2/X vssd1 vssd1 vccd1 vccd1 _6360_/X sky130_fd_sc_hd__or2_1
X_5311_ _5605_/B vssd1 vssd1 vccd1 vccd1 _6966_/A sky130_fd_sc_hd__clkbuf_4
X_6291_ _6528_/B _6290_/B _6290_/C vssd1 vssd1 vccd1 vccd1 _6292_/B sky130_fd_sc_hd__a21oi_1
X_5242_ _5242_/A _5242_/B vssd1 vssd1 vccd1 vccd1 _5245_/A sky130_fd_sc_hd__xnor2_4
X_5173_ _5173_/A _5173_/B vssd1 vssd1 vccd1 vccd1 _5176_/A sky130_fd_sc_hd__nand2_2
X_4124_ _4124_/A vssd1 vssd1 vccd1 vccd1 _4375_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput1 active vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_4
XFILLER_83_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4055_ _7162_/Q vssd1 vssd1 vccd1 vccd1 _4795_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_71_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4957_ _4957_/A _5121_/A _4957_/C vssd1 vssd1 vccd1 vccd1 _5277_/B sky130_fd_sc_hd__and3_1
X_4888_ _4888_/A _4888_/B vssd1 vssd1 vccd1 vccd1 _4907_/A sky130_fd_sc_hd__xor2_1
X_3908_ _3908_/A _3908_/B vssd1 vssd1 vccd1 vccd1 _3909_/B sky130_fd_sc_hd__xor2_1
X_3839_ _4613_/A _5125_/A _3838_/Y vssd1 vssd1 vccd1 vccd1 _4011_/A sky130_fd_sc_hd__a21o_2
X_6627_ _6627_/A vssd1 vssd1 vccd1 vccd1 _6973_/A sky130_fd_sc_hd__inv_2
X_6558_ _6718_/A _6718_/B vssd1 vssd1 vccd1 vccd1 _6583_/A sky130_fd_sc_hd__xor2_1
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6489_ _6491_/A _6491_/B _6492_/B vssd1 vssd1 vccd1 vccd1 _6514_/B sky130_fd_sc_hd__and3_1
X_5509_ _5510_/A _5510_/B _5510_/C vssd1 vssd1 vccd1 vccd1 _5558_/A sky130_fd_sc_hd__o21ai_1
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5860_ _5860_/A _5860_/B vssd1 vssd1 vccd1 vccd1 _5861_/B sky130_fd_sc_hd__nor2_2
X_4811_ _4865_/A _4813_/B _4810_/X vssd1 vssd1 vccd1 vccd1 _4931_/A sky130_fd_sc_hd__o21ai_1
XFILLER_61_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5791_ _5792_/A _5792_/B vssd1 vssd1 vccd1 vccd1 _6076_/A sky130_fd_sc_hd__and2_1
X_4742_ _4742_/A _4742_/B vssd1 vssd1 vccd1 vccd1 _4748_/A sky130_fd_sc_hd__xor2_1
X_4673_ _5872_/A vssd1 vssd1 vccd1 vccd1 _6137_/B sky130_fd_sc_hd__buf_4
X_3624_ _3648_/A vssd1 vssd1 vccd1 vccd1 _3629_/A sky130_fd_sc_hd__buf_8
X_6412_ _6586_/B _6586_/A vssd1 vssd1 vccd1 vccd1 _6607_/B sky130_fd_sc_hd__or2b_1
X_7392_ _7392_/A _3684_/Y vssd1 vssd1 vccd1 vccd1 io_out[34] sky130_fd_sc_hd__ebufn_8
X_6343_ _6297_/A _6297_/B _6342_/X vssd1 vssd1 vccd1 vccd1 _6380_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6274_ _6274_/A _6274_/B _6274_/C vssd1 vssd1 vccd1 vccd1 _6324_/C sky130_fd_sc_hd__nand3_1
XFILLER_88_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5225_ _5690_/A _5719_/A vssd1 vssd1 vccd1 vccd1 _5226_/B sky130_fd_sc_hd__nor2_1
XFILLER_69_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5156_ _5156_/A _5033_/B vssd1 vssd1 vccd1 vccd1 _5156_/X sky130_fd_sc_hd__or2b_1
XFILLER_96_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4107_ _7164_/Q vssd1 vssd1 vccd1 vccd1 _5021_/A sky130_fd_sc_hd__buf_2
XFILLER_56_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5087_ _5236_/B _5087_/B vssd1 vssd1 vccd1 vccd1 _5088_/B sky130_fd_sc_hd__xnor2_2
X_4038_ _4038_/A _4038_/B vssd1 vssd1 vccd1 vccd1 _4187_/B sky130_fd_sc_hd__nor2_4
XFILLER_37_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5989_ _5989_/A _5989_/B vssd1 vssd1 vccd1 vccd1 _5990_/B sky130_fd_sc_hd__nand2_1
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_50 _7117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7259__52 vssd1 vssd1 vccd1 vccd1 _7259__52/HI _7358_/A sky130_fd_sc_hd__conb_1
XFILLER_97_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_3_4_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7172_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _5719_/A vssd1 vssd1 vccd1 vccd1 _6140_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_97_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6961_ _6475_/A _6949_/X _6960_/X _6952_/X vssd1 vssd1 vccd1 vccd1 _7164_/D sky130_fd_sc_hd__o211a_1
XFILLER_19_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5912_ _5912_/A _5912_/B vssd1 vssd1 vccd1 vccd1 _5913_/B sky130_fd_sc_hd__nand2_1
X_6892_ _6893_/B vssd1 vssd1 vccd1 vccd1 _6892_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5843_ _5775_/Y _5823_/X _5841_/B _5842_/Y vssd1 vssd1 vccd1 vccd1 _5844_/B sky130_fd_sc_hd__a31oi_4
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5774_ _5774_/A _5774_/B vssd1 vssd1 vccd1 vccd1 _5840_/B sky130_fd_sc_hd__xnor2_1
X_4725_ _6933_/A _4803_/B vssd1 vssd1 vccd1 vccd1 _4759_/A sky130_fd_sc_hd__or2_1
X_4656_ _4656_/A _4656_/B vssd1 vssd1 vccd1 vccd1 _4691_/A sky130_fd_sc_hd__nor2_1
X_7375_ _7375_/A _3664_/Y vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__ebufn_8
X_4587_ _4587_/A _4587_/B vssd1 vssd1 vccd1 vccd1 _4663_/A sky130_fd_sc_hd__xnor2_1
X_6326_ _6264_/A _6268_/Y _6270_/X vssd1 vssd1 vccd1 vccd1 _6327_/B sky130_fd_sc_hd__a21bo_1
XFILLER_88_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6257_ _6258_/A _6258_/B vssd1 vssd1 vccd1 vccd1 _6257_/X sky130_fd_sc_hd__or2_1
XFILLER_57_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6188_ _6188_/A _6252_/B vssd1 vssd1 vccd1 vccd1 _6255_/A sky130_fd_sc_hd__xor2_4
X_5208_ _5335_/A _5208_/B vssd1 vssd1 vccd1 vccd1 _5210_/A sky130_fd_sc_hd__nor2_1
XFILLER_29_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5139_ _5266_/A _5139_/B vssd1 vssd1 vccd1 vccd1 _5141_/C sky130_fd_sc_hd__xnor2_1
XFILLER_84_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7307__100 vssd1 vssd1 vccd1 vccd1 _7307__100/HI _7415_/A sky130_fd_sc_hd__conb_1
X_4510_ _4511_/A _4511_/B vssd1 vssd1 vccd1 vccd1 _4607_/B sky130_fd_sc_hd__xor2_2
X_5490_ _5490_/A _5490_/B _5490_/C vssd1 vssd1 vccd1 vccd1 _5491_/B sky130_fd_sc_hd__or3_1
X_4441_ _4439_/A _4439_/B _4493_/A vssd1 vssd1 vccd1 vccd1 _4444_/A sky130_fd_sc_hd__a21o_1
Xhold106 _4856_/A vssd1 vssd1 vccd1 vccd1 _7102_/A sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold117 hold25/X vssd1 vssd1 vccd1 vccd1 hold117/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_7160_ _7225_/CLK _7160_/D vssd1 vssd1 vccd1 vccd1 _7160_/Q sky130_fd_sc_hd__dfxtp_1
Xhold128 hold41/X vssd1 vssd1 vccd1 vccd1 hold128/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_6111_ _6111_/A _6111_/B vssd1 vssd1 vccd1 vccd1 _6112_/A sky130_fd_sc_hd__nand2_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4372_ _4372_/A _4372_/B vssd1 vssd1 vccd1 vccd1 _4382_/A sky130_fd_sc_hd__nor2_1
XFILLER_98_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7091_ _7091_/A _7091_/B vssd1 vssd1 vccd1 vccd1 _7091_/X sky130_fd_sc_hd__or2_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6042_ _6142_/B _6999_/A vssd1 vssd1 vccd1 vccd1 _6047_/A sky130_fd_sc_hd__nand2_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6944_ input7/X _6935_/X _6943_/X _6939_/X vssd1 vssd1 vccd1 vccd1 _7158_/D sky130_fd_sc_hd__o211a_1
XFILLER_81_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6875_ _6875_/A _6875_/B vssd1 vssd1 vccd1 vccd1 _6876_/B sky130_fd_sc_hd__nand2_1
XFILLER_22_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5826_ _5826_/A _5826_/B vssd1 vssd1 vccd1 vccd1 _5836_/B sky130_fd_sc_hd__xor2_1
XFILLER_22_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5757_ _5756_/Y _5897_/B _5628_/Y vssd1 vssd1 vccd1 vccd1 _5838_/B sky130_fd_sc_hd__a21oi_2
X_4708_ _4707_/A _4708_/B vssd1 vssd1 vccd1 vccd1 _4708_/X sky130_fd_sc_hd__and2b_1
X_7427_ _7427_/A _3725_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[31] sky130_fd_sc_hd__ebufn_8
X_5688_ _5688_/A _5688_/B vssd1 vssd1 vccd1 vccd1 _6049_/A sky130_fd_sc_hd__xor2_4
X_4639_ _7078_/A _4639_/B vssd1 vssd1 vccd1 vccd1 _4695_/B sky130_fd_sc_hd__xnor2_1
X_7358_ _7358_/A _3736_/Y vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__ebufn_8
XFILLER_78_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6309_ _6309_/A _6354_/A vssd1 vssd1 vccd1 vccd1 _6313_/A sky130_fd_sc_hd__xnor2_2
X_7229__22 vssd1 vssd1 vccd1 vccd1 _7229__22/HI _7328_/A sky130_fd_sc_hd__conb_1
XFILLER_94_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4990_ _5287_/A _4990_/B vssd1 vssd1 vccd1 vccd1 _4992_/C sky130_fd_sc_hd__xnor2_1
X_3941_ _4799_/A _5121_/A vssd1 vssd1 vccd1 vccd1 _3978_/B sky130_fd_sc_hd__nor2_1
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3872_ _3908_/A _3978_/A _3907_/B _3867_/B _3867_/A vssd1 vssd1 vccd1 vccd1 _4981_/A
+ sky130_fd_sc_hd__o32a_1
X_6660_ _6659_/Y _6679_/B _3781_/X vssd1 vssd1 vccd1 vccd1 _6662_/B sky130_fd_sc_hd__o21ai_1
XFILLER_31_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5611_ _6571_/A _6589_/A _5611_/C vssd1 vssd1 vccd1 vccd1 _5636_/A sky130_fd_sc_hd__and3_1
X_6591_ _6978_/A _6589_/B _6622_/A vssd1 vssd1 vccd1 vccd1 _6594_/B sky130_fd_sc_hd__o21ai_2
X_5542_ _5542_/A _5542_/B vssd1 vssd1 vccd1 vccd1 _5543_/B sky130_fd_sc_hd__xnor2_1
X_5473_ _5531_/B _5472_/Y hold63/X vssd1 vssd1 vccd1 vccd1 _5473_/X sky130_fd_sc_hd__a21o_1
X_4424_ _7153_/Q vssd1 vssd1 vccd1 vccd1 _6502_/B sky130_fd_sc_hd__buf_2
X_7212_ _7222_/CLK hold88/X vssd1 vssd1 vccd1 vccd1 _7212_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_98_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4355_ _4355_/A _5056_/C vssd1 vssd1 vccd1 vccd1 _4363_/A sky130_fd_sc_hd__or2_1
X_7143_ _7226_/CLK hold24/X vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__dfxtp_1
X_7074_ hold119/X _7062_/X _7072_/Y _7073_/X vssd1 vssd1 vccd1 vccd1 _7206_/D sky130_fd_sc_hd__o211a_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4286_ _4286_/A vssd1 vssd1 vccd1 vccd1 _6045_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_100_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6025_ _6107_/A _6107_/B vssd1 vssd1 vccd1 vccd1 _6033_/A sky130_fd_sc_hd__xnor2_4
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6927_ input18/X _7116_/B _6926_/X _6846_/X vssd1 vssd1 vccd1 vccd1 _7152_/D sky130_fd_sc_hd__o211a_1
X_6858_ _6859_/A _6859_/B vssd1 vssd1 vccd1 vccd1 _6875_/A sky130_fd_sc_hd__nand2_1
XFILLER_50_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5809_ _5434_/B _5802_/B _5815_/B _5815_/A vssd1 vssd1 vccd1 vccd1 _6084_/A sky130_fd_sc_hd__o2bb2a_2
X_6789_ _6789_/A _6789_/B vssd1 vssd1 vccd1 vccd1 _6789_/Y sky130_fd_sc_hd__nand2_2
XFILLER_13_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4140_ _4279_/A _5002_/A vssd1 vssd1 vccd1 vccd1 _5006_/B sky130_fd_sc_hd__and2b_1
X_4071_ _4215_/A _4215_/B vssd1 vssd1 vccd1 vccd1 _4216_/A sky130_fd_sc_hd__nand2_1
XFILLER_83_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4973_ _4974_/A _4974_/B vssd1 vssd1 vccd1 vccd1 _4975_/A sky130_fd_sc_hd__or2_1
XFILLER_36_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3924_ _5671_/B vssd1 vssd1 vccd1 vccd1 _4506_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_6712_ _6679_/A _6421_/A _6420_/B _6423_/Y vssd1 vssd1 vccd1 vccd1 _6715_/B sky130_fd_sc_hd__o31a_1
XFILLER_51_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6643_ _6643_/A _6643_/B vssd1 vssd1 vccd1 vccd1 _6644_/B sky130_fd_sc_hd__xnor2_1
X_3855_ _3877_/C _3896_/A vssd1 vssd1 vccd1 vccd1 _3920_/A sky130_fd_sc_hd__xor2_2
X_6574_ _6736_/A _6596_/B _6573_/Y vssd1 vssd1 vccd1 vccd1 _6576_/A sky130_fd_sc_hd__a21o_1
X_3786_ _3785_/B _3785_/C _3785_/A vssd1 vssd1 vccd1 vccd1 _3787_/B sky130_fd_sc_hd__a21oi_1
X_5525_ _5525_/A _5525_/B vssd1 vssd1 vccd1 vccd1 _5526_/B sky130_fd_sc_hd__nor2_1
X_5456_ _5456_/A _5456_/B vssd1 vssd1 vccd1 vccd1 _5518_/A sky130_fd_sc_hd__xnor2_1
X_4407_ _4407_/A _4407_/B _4407_/C vssd1 vssd1 vccd1 vccd1 _4407_/X sky130_fd_sc_hd__or3_1
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5387_ _5387_/A _5387_/B vssd1 vssd1 vccd1 vccd1 _5399_/A sky130_fd_sc_hd__nor2_1
XFILLER_86_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4338_ _4338_/A _4338_/B vssd1 vssd1 vccd1 vccd1 _4442_/A sky130_fd_sc_hd__xor2_1
X_7126_ _7226_/CLK hold62/X vssd1 vssd1 vccd1 vccd1 hold61/A sky130_fd_sc_hd__dfxtp_1
XFILLER_75_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7057_ hold97/X _7059_/B vssd1 vssd1 vccd1 vccd1 _7057_/X sky130_fd_sc_hd__or2_1
XFILLER_47_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4269_ _4317_/A vssd1 vssd1 vccd1 vccd1 _4466_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_101_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6008_ _6007_/A _5967_/Y _5935_/Y vssd1 vssd1 vccd1 vccd1 _6009_/C sky130_fd_sc_hd__o21ai_1
XFILLER_55_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3640_ _3641_/A vssd1 vssd1 vccd1 vccd1 _3640_/Y sky130_fd_sc_hd__inv_2
X_5310_ _5606_/B vssd1 vssd1 vccd1 vccd1 _5605_/B sky130_fd_sc_hd__inv_2
X_6290_ _6528_/B _6290_/B _6290_/C vssd1 vssd1 vccd1 vccd1 _6346_/B sky130_fd_sc_hd__and3_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5241_ _5365_/B _5241_/B vssd1 vssd1 vccd1 vccd1 _5242_/B sky130_fd_sc_hd__xor2_4
XFILLER_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5172_ _5171_/A _5171_/B _5171_/C vssd1 vssd1 vccd1 vccd1 _5173_/B sky130_fd_sc_hd__a21o_1
XFILLER_29_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4123_ _5011_/A _7180_/Q vssd1 vssd1 vccd1 vccd1 _4124_/A sky130_fd_sc_hd__and2_1
Xinput2 io_in[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4054_ _4054_/A _4078_/A vssd1 vssd1 vccd1 vccd1 _4065_/A sky130_fd_sc_hd__or2_1
XFILLER_68_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4956_ _7214_/Q _4956_/B vssd1 vssd1 vccd1 vccd1 _4957_/C sky130_fd_sc_hd__or2_1
X_4887_ _4925_/B _4887_/B vssd1 vssd1 vccd1 vccd1 _4888_/B sky130_fd_sc_hd__xnor2_1
X_3907_ _3978_/A _3907_/B vssd1 vssd1 vccd1 vccd1 _3908_/B sky130_fd_sc_hd__or2_1
XFILLER_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3838_ _6027_/A _5722_/A vssd1 vssd1 vccd1 vccd1 _3838_/Y sky130_fd_sc_hd__nor2_1
X_6626_ _6627_/A _6624_/X _6657_/A vssd1 vssd1 vccd1 vccd1 _6628_/B sky130_fd_sc_hd__a21oi_1
X_6557_ _6717_/A _6717_/B vssd1 vssd1 vccd1 vccd1 _6718_/B sky130_fd_sc_hd__xnor2_1
X_3769_ _4356_/B _3807_/A vssd1 vssd1 vccd1 vccd1 _3801_/B sky130_fd_sc_hd__xnor2_1
X_5508_ _5508_/A _5508_/B vssd1 vssd1 vccd1 vccd1 _5510_/C sky130_fd_sc_hd__xnor2_1
X_6488_ _6110_/A _6466_/A _6466_/B _6487_/X vssd1 vssd1 vccd1 vccd1 _6492_/B sky130_fd_sc_hd__a31o_1
X_5439_ _5216_/A _5337_/B hold82/A vssd1 vssd1 vccd1 vccd1 _5547_/B sky130_fd_sc_hd__a21oi_2
XFILLER_101_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7109_ _5292_/A _7101_/X _7108_/X _7099_/X vssd1 vssd1 vccd1 vccd1 _7109_/X sky130_fd_sc_hd__o211a_1
XFILLER_59_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4810_ _4810_/A _4809_/A vssd1 vssd1 vccd1 vccd1 _4810_/X sky130_fd_sc_hd__or2b_1
XFILLER_33_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5790_ _5435_/A _5802_/A _5434_/Y vssd1 vssd1 vccd1 vccd1 _5792_/B sky130_fd_sc_hd__o21a_1
X_4741_ _4741_/A _4741_/B vssd1 vssd1 vccd1 vccd1 _4742_/A sky130_fd_sc_hd__xnor2_1
X_4672_ _4676_/A _4741_/B vssd1 vssd1 vccd1 vccd1 _4672_/Y sky130_fd_sc_hd__nor2_1
X_3623_ input1/X vssd1 vssd1 vccd1 vccd1 _3648_/A sky130_fd_sc_hd__clkbuf_4
X_6411_ _6560_/A _6411_/B vssd1 vssd1 vccd1 vccd1 _6586_/A sky130_fd_sc_hd__xnor2_2
X_7391_ _7391_/A _3683_/Y vssd1 vssd1 vccd1 vccd1 io_out[33] sky130_fd_sc_hd__ebufn_8
X_6342_ _6342_/A _6285_/A vssd1 vssd1 vccd1 vccd1 _6342_/X sky130_fd_sc_hd__or2b_1
X_6273_ _6274_/A _6274_/B _6274_/C vssd1 vssd1 vccd1 vccd1 _6327_/A sky130_fd_sc_hd__a21o_1
X_5224_ _6034_/A vssd1 vssd1 vccd1 vccd1 _6129_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5155_ _5321_/A _5155_/B vssd1 vssd1 vccd1 vccd1 _5265_/A sky130_fd_sc_hd__and2b_1
XFILLER_84_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4106_ _7165_/Q vssd1 vssd1 vccd1 vccd1 _4279_/A sky130_fd_sc_hd__clkbuf_2
X_5086_ _5086_/A _5086_/B vssd1 vssd1 vccd1 vccd1 _5087_/B sky130_fd_sc_hd__or2_1
X_4037_ _4036_/A _4036_/B _4036_/C vssd1 vssd1 vccd1 vccd1 _4038_/B sky130_fd_sc_hd__a21oi_1
XFILLER_56_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5988_ _5989_/A _5989_/B vssd1 vssd1 vccd1 vccd1 _5990_/A sky130_fd_sc_hd__or2_1
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4939_ _4836_/A _4838_/X _4787_/Y vssd1 vssd1 vccd1 vccd1 _4939_/Y sky130_fd_sc_hd__o21bai_2
XANTENNA_40 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_51 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6609_ _6609_/A _6609_/B vssd1 vssd1 vccd1 vccd1 _6609_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7324__117 vssd1 vssd1 vccd1 vccd1 _7324__117/HI _7432_/A sky130_fd_sc_hd__conb_1
XFILLER_97_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7274__67 vssd1 vssd1 vccd1 vccd1 _7274__67/HI _7373_/A sky130_fd_sc_hd__conb_1
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6960_ _6960_/A _6975_/B vssd1 vssd1 vccd1 vccd1 _6960_/X sky130_fd_sc_hd__or2_1
X_5911_ _5911_/A _5911_/B vssd1 vssd1 vccd1 vccd1 _5948_/A sky130_fd_sc_hd__xor2_4
XFILLER_19_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6891_ input9/X _6891_/B _6891_/C vssd1 vssd1 vccd1 vccd1 _6893_/B sky130_fd_sc_hd__and3b_4
X_5842_ _5868_/A _5868_/B vssd1 vssd1 vccd1 vccd1 _5842_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5773_ _5773_/A _5773_/B vssd1 vssd1 vccd1 vccd1 _5840_/A sky130_fd_sc_hd__nor2_1
XFILLER_61_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4724_ _4741_/A _4724_/B vssd1 vssd1 vccd1 vccd1 _4803_/B sky130_fd_sc_hd__nand2_1
X_4655_ _4655_/A _4703_/A _4655_/C vssd1 vssd1 vccd1 vccd1 _4656_/B sky130_fd_sc_hd__and3_1
X_4586_ _4586_/A _4586_/B vssd1 vssd1 vccd1 vccd1 _4587_/A sky130_fd_sc_hd__or2_1
X_7374_ _7374_/A _3663_/Y vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__ebufn_8
X_6325_ _6325_/A _6325_/B vssd1 vssd1 vccd1 vccd1 _6332_/B sky130_fd_sc_hd__nor2_1
XFILLER_67_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6256_ _6194_/A _6194_/B _6255_/X vssd1 vssd1 vccd1 vccd1 _6258_/B sky130_fd_sc_hd__o21ai_2
X_5207_ hold82/A hold87/A hold53/A vssd1 vssd1 vccd1 vccd1 _5208_/B sky130_fd_sc_hd__a21oi_1
X_6187_ _6089_/A _6089_/B _6186_/X vssd1 vssd1 vccd1 vccd1 _6252_/B sky130_fd_sc_hd__o21ai_4
XFILLER_84_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5138_ _5266_/B _5289_/B vssd1 vssd1 vccd1 vccd1 _5139_/B sky130_fd_sc_hd__nand2_1
XFILLER_83_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5069_ _5341_/A _5341_/B vssd1 vssd1 vccd1 vccd1 _5220_/B sky130_fd_sc_hd__xnor2_1
XFILLER_80_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4440_ _4492_/B _4440_/B vssd1 vssd1 vccd1 vccd1 _4493_/A sky130_fd_sc_hd__and2b_1
Xhold107 _7103_/X vssd1 vssd1 vccd1 vccd1 _7217_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold118 hold30/X vssd1 vssd1 vccd1 vccd1 hold118/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_6110_ _6110_/A _6109_/A vssd1 vssd1 vccd1 vccd1 _6111_/B sky130_fd_sc_hd__or2b_1
X_4371_ _4301_/A _4301_/B _4370_/Y vssd1 vssd1 vccd1 vccd1 _4384_/A sky130_fd_sc_hd__a21bo_1
X_7090_ hold87/X _7088_/X _7089_/Y _7086_/X vssd1 vssd1 vccd1 vccd1 hold88/A sky130_fd_sc_hd__o211a_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6041_ _6147_/B _6041_/B vssd1 vssd1 vccd1 vccd1 _6048_/A sky130_fd_sc_hd__xor2_4
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6943_ _6943_/A _6954_/B vssd1 vssd1 vccd1 vccd1 _6943_/X sky130_fd_sc_hd__or2_1
XFILLER_54_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6874_ _6874_/A _6874_/B vssd1 vssd1 vccd1 vccd1 _6876_/A sky130_fd_sc_hd__xor2_1
X_5825_ _6999_/A _6997_/A vssd1 vssd1 vccd1 vccd1 _5870_/A sky130_fd_sc_hd__and2_1
X_5756_ _5756_/A vssd1 vssd1 vccd1 vccd1 _5756_/Y sky130_fd_sc_hd__inv_2
X_4707_ _4707_/A _4708_/B vssd1 vssd1 vccd1 vccd1 _4758_/B sky130_fd_sc_hd__xnor2_2
X_5687_ _5687_/A _5687_/B vssd1 vssd1 vccd1 vccd1 _5688_/B sky130_fd_sc_hd__xnor2_2
X_7426_ _7426_/A _3724_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[30] sky130_fd_sc_hd__ebufn_8
X_4638_ _7038_/A _4638_/B vssd1 vssd1 vccd1 vccd1 _4695_/A sky130_fd_sc_hd__nand2_1
X_7357_ _7357_/A _3645_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[31] sky130_fd_sc_hd__ebufn_8
XFILLER_89_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4569_ _4569_/A _4569_/B vssd1 vssd1 vccd1 vccd1 _4570_/B sky130_fd_sc_hd__xnor2_1
X_6308_ _6306_/Y _6246_/B _6307_/Y vssd1 vssd1 vccd1 vccd1 _6354_/A sky130_fd_sc_hd__a21oi_1
X_6239_ _6166_/A _6166_/B _6169_/B vssd1 vssd1 vccd1 vccd1 _6244_/A sky130_fd_sc_hd__a21o_1
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7244__37 vssd1 vssd1 vccd1 vccd1 _7244__37/HI _7343_/A sky130_fd_sc_hd__conb_1
XFILLER_84_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3940_ _7214_/Q _4956_/B vssd1 vssd1 vccd1 vccd1 _5121_/A sky130_fd_sc_hd__nand2_1
XFILLER_44_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3871_ _5131_/A _7083_/A vssd1 vssd1 vccd1 vccd1 _3907_/B sky130_fd_sc_hd__nor2_1
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6590_ _6625_/A _6621_/B vssd1 vssd1 vccd1 vccd1 _6622_/A sky130_fd_sc_hd__nand2_1
X_5610_ _5737_/A vssd1 vssd1 vccd1 vccd1 _6589_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5541_ _7055_/A _5541_/B vssd1 vssd1 vccd1 vccd1 _5542_/A sky130_fd_sc_hd__or2_1
X_7211_ _7221_/CLK _7211_/D vssd1 vssd1 vccd1 vccd1 _7211_/Q sky130_fd_sc_hd__dfxtp_1
X_5472_ _5472_/A _5472_/B _5472_/C vssd1 vssd1 vccd1 vccd1 _5472_/Y sky130_fd_sc_hd__nand3_1
X_4423_ _4553_/A vssd1 vssd1 vccd1 vccd1 _6475_/A sky130_fd_sc_hd__clkbuf_4
X_7142_ _7224_/CLK _7142_/D vssd1 vssd1 vccd1 vccd1 hold65/A sky130_fd_sc_hd__dfxtp_1
X_4354_ _4354_/A vssd1 vssd1 vccd1 vccd1 _5056_/C sky130_fd_sc_hd__inv_2
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7073_ _7073_/A vssd1 vssd1 vccd1 vccd1 _7073_/X sky130_fd_sc_hd__clkbuf_2
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6024_ _6106_/A _6106_/B _6021_/X _6023_/Y vssd1 vssd1 vccd1 vccd1 _6107_/B sky130_fd_sc_hd__a211o_2
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4285_ _4285_/A _4285_/B vssd1 vssd1 vccd1 vccd1 _4289_/A sky130_fd_sc_hd__nor2_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6926_ _6926_/A _6954_/B vssd1 vssd1 vccd1 vccd1 _6926_/X sky130_fd_sc_hd__or2_1
XFILLER_54_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6857_ _6828_/A _6828_/B _6856_/X vssd1 vssd1 vccd1 vccd1 _6859_/B sky130_fd_sc_hd__a21bo_1
X_6788_ _6789_/A _6789_/B vssd1 vssd1 vccd1 vccd1 _6788_/X sky130_fd_sc_hd__or2_1
X_5808_ _5854_/A _5808_/B vssd1 vssd1 vccd1 vccd1 _5815_/A sky130_fd_sc_hd__xnor2_2
XFILLER_50_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5739_ _5745_/A _5736_/X _5787_/B _5739_/D vssd1 vssd1 vccd1 vccd1 _5745_/B sky130_fd_sc_hd__and4bb_1
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7409_ _7409_/A _3705_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[13] sky130_fd_sc_hd__ebufn_8
XFILLER_89_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4070_ _4070_/A _4070_/B vssd1 vssd1 vccd1 vccd1 _4215_/B sky130_fd_sc_hd__nor2_1
XFILLER_95_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4972_ _4972_/A _5145_/C vssd1 vssd1 vccd1 vccd1 _4974_/B sky130_fd_sc_hd__xnor2_1
X_3923_ _7185_/Q _7184_/Q vssd1 vssd1 vccd1 vccd1 _5671_/B sky130_fd_sc_hd__xor2_4
X_6711_ _6711_/A _6711_/B vssd1 vssd1 vccd1 vccd1 _6750_/B sky130_fd_sc_hd__nand2_1
XFILLER_32_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3854_ _4003_/A _7198_/Q vssd1 vssd1 vccd1 vccd1 _3896_/A sky130_fd_sc_hd__nand2_1
X_6642_ _6650_/A _6650_/B _6641_/X vssd1 vssd1 vccd1 vccd1 _6645_/B sky130_fd_sc_hd__a21o_1
X_6573_ _6573_/A _6573_/B vssd1 vssd1 vccd1 vccd1 _6573_/Y sky130_fd_sc_hd__nor2_1
X_3785_ _3785_/A _3785_/B _3785_/C vssd1 vssd1 vccd1 vccd1 _4353_/A sky130_fd_sc_hd__and3_2
X_5524_ _5524_/A _5524_/B vssd1 vssd1 vccd1 vccd1 _5525_/B sky130_fd_sc_hd__and2_1
X_5455_ _5499_/A _5499_/B vssd1 vssd1 vccd1 vccd1 _5456_/B sky130_fd_sc_hd__xor2_1
X_4406_ _4406_/A _4406_/B vssd1 vssd1 vccd1 vccd1 _4407_/C sky130_fd_sc_hd__and2_1
XFILLER_99_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7125_ _7226_/CLK hold57/X vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__dfxtp_1
X_5386_ _5386_/A _5386_/B _5386_/C vssd1 vssd1 vccd1 vccd1 _5387_/B sky130_fd_sc_hd__nor3_1
X_4337_ _4445_/A _4445_/B _4336_/X vssd1 vssd1 vccd1 vccd1 _4338_/B sky130_fd_sc_hd__a21oi_2
XFILLER_86_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7056_ hold125/X _7045_/X _7055_/Y _7048_/X vssd1 vssd1 vccd1 vccd1 _7199_/D sky130_fd_sc_hd__o211a_1
X_4268_ _7182_/Q _4377_/B vssd1 vssd1 vccd1 vccd1 _4272_/A sky130_fd_sc_hd__xnor2_1
XFILLER_101_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6007_ _6007_/A _6007_/B vssd1 vssd1 vccd1 vccd1 _6009_/B sky130_fd_sc_hd__nand2_1
X_4199_ _4195_/A _4194_/A _4416_/B _4406_/A vssd1 vssd1 vccd1 vccd1 _4238_/B sky130_fd_sc_hd__o31a_1
XFILLER_39_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6909_ hold10/X _6890_/X _6908_/X vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__a21oi_1
XFILLER_23_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5240_ _5364_/B _5240_/B vssd1 vssd1 vccd1 vccd1 _5241_/B sky130_fd_sc_hd__xor2_2
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5171_ _5171_/A _5171_/B _5171_/C vssd1 vssd1 vccd1 vccd1 _5173_/A sky130_fd_sc_hd__nand3_1
X_4122_ _7181_/Q vssd1 vssd1 vccd1 vccd1 _5011_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4053_ _4054_/A _4053_/B _4070_/A vssd1 vssd1 vccd1 vccd1 _4078_/A sky130_fd_sc_hd__nor3b_1
XFILLER_68_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput3 io_in[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_2
XFILLER_49_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4955_ _5127_/A _4955_/B vssd1 vssd1 vccd1 vccd1 _5119_/A sky130_fd_sc_hd__nor2_1
XFILLER_51_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3906_ _3921_/A _3921_/B _3905_/Y vssd1 vssd1 vccd1 vccd1 _3965_/A sky130_fd_sc_hd__o21ba_1
XFILLER_51_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4886_ _4886_/A _4890_/A vssd1 vssd1 vccd1 vccd1 _4887_/B sky130_fd_sc_hd__nor2_1
X_3837_ _7187_/Q vssd1 vssd1 vccd1 vccd1 _5722_/A sky130_fd_sc_hd__clkbuf_2
X_6625_ _6625_/A _6625_/B vssd1 vssd1 vccd1 vccd1 _6657_/A sky130_fd_sc_hd__and2_1
X_3768_ _7066_/A hold98/A vssd1 vssd1 vccd1 vccd1 _3807_/A sky130_fd_sc_hd__and2_1
XFILLER_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6556_ _6579_/A _6579_/B _6555_/X vssd1 vssd1 vccd1 vccd1 _6717_/B sky130_fd_sc_hd__a21oi_2
X_5507_ _5507_/A _5507_/B vssd1 vssd1 vccd1 vccd1 _5508_/B sky130_fd_sc_hd__nand2_1
X_6487_ _6487_/A _6487_/B _6487_/C _6487_/D vssd1 vssd1 vccd1 vccd1 _6487_/X sky130_fd_sc_hd__and4_1
X_3699_ _3703_/A vssd1 vssd1 vccd1 vccd1 _3699_/Y sky130_fd_sc_hd__inv_2
X_5438_ _5438_/A vssd1 vssd1 vccd1 vccd1 _5547_/A sky130_fd_sc_hd__inv_2
X_5369_ _5249_/A _5249_/B _5368_/X vssd1 vssd1 vccd1 vccd1 _5468_/B sky130_fd_sc_hd__a21oi_2
X_7108_ _7108_/A _7114_/B vssd1 vssd1 vccd1 vccd1 _7108_/X sky130_fd_sc_hd__or2_1
XFILLER_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7039_ hold111/X _7032_/X _7038_/X _7034_/X vssd1 vssd1 vccd1 vccd1 _7193_/D sky130_fd_sc_hd__o211a_1
XFILLER_47_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4740_ _4754_/A _4754_/B vssd1 vssd1 vccd1 vccd1 _4757_/A sky130_fd_sc_hd__xnor2_1
XFILLER_61_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4671_ _4671_/A _4671_/B vssd1 vssd1 vccd1 vccd1 _4741_/B sky130_fd_sc_hd__and2_1
X_3622_ _3622_/A vssd1 vssd1 vccd1 vccd1 _3622_/Y sky130_fd_sc_hd__inv_2
X_7390_ _7390_/A _3682_/Y vssd1 vssd1 vccd1 vccd1 io_out[32] sky130_fd_sc_hd__ebufn_8
X_6410_ _6410_/A _6559_/A vssd1 vssd1 vccd1 vccd1 _6411_/B sky130_fd_sc_hd__xnor2_1
X_6341_ _6341_/A _6341_/B vssd1 vssd1 vccd1 vccd1 _6344_/A sky130_fd_sc_hd__xnor2_1
X_6272_ _5450_/B _6268_/Y _6270_/X _6271_/Y vssd1 vssd1 vccd1 vccd1 _6274_/C sky130_fd_sc_hd__a22oi_1
X_5223_ _5218_/A _4267_/B _5083_/B _5086_/B vssd1 vssd1 vccd1 vccd1 _5354_/B sky130_fd_sc_hd__a31o_1
XFILLER_69_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5154_ _5154_/A _5154_/B vssd1 vssd1 vccd1 vccd1 _5155_/B sky130_fd_sc_hd__or2_1
X_4105_ _4372_/A _4372_/B vssd1 vssd1 vccd1 vccd1 _4117_/A sky130_fd_sc_hd__xnor2_1
X_5085_ _5689_/A _5085_/B vssd1 vssd1 vccd1 vccd1 _5086_/B sky130_fd_sc_hd__and2_1
X_4036_ _4036_/A _4036_/B _4036_/C vssd1 vssd1 vccd1 vccd1 _4038_/A sky130_fd_sc_hd__and3_1
XFILLER_71_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5987_ _5987_/A _6577_/A _5987_/C vssd1 vssd1 vccd1 vccd1 _5989_/B sky130_fd_sc_hd__and3_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4938_ _4940_/A _4940_/B vssd1 vssd1 vccd1 vccd1 _4938_/X sky130_fd_sc_hd__or2_1
XFILLER_12_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4869_ _4869_/A _4869_/B vssd1 vssd1 vccd1 vccd1 _4925_/B sky130_fd_sc_hd__xor2_1
XANTENNA_30 _3672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_41 _6627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_52 _7007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6608_ _6711_/A _6608_/B vssd1 vssd1 vccd1 vccd1 _6643_/B sky130_fd_sc_hd__or2_1
X_6539_ _6539_/A _6539_/B vssd1 vssd1 vccd1 vccd1 _6540_/B sky130_fd_sc_hd__and2_1
XFILLER_97_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5910_ _5910_/A _5910_/B vssd1 vssd1 vccd1 vccd1 _5918_/A sky130_fd_sc_hd__or2_1
X_6890_ _6893_/A vssd1 vssd1 vccd1 vccd1 _6890_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5841_ _5841_/A _5841_/B vssd1 vssd1 vccd1 vccd1 _5868_/B sky130_fd_sc_hd__xor2_1
X_5772_ _5714_/A _4852_/Y _5750_/B vssd1 vssd1 vccd1 vccd1 _5773_/B sky130_fd_sc_hd__a21boi_1
X_4723_ _4723_/A _4723_/B vssd1 vssd1 vccd1 vccd1 _4724_/B sky130_fd_sc_hd__or2_1
X_4654_ _4655_/A _4703_/A _4655_/C vssd1 vssd1 vccd1 vccd1 _4656_/A sky130_fd_sc_hd__a21oi_1
X_4585_ _4658_/A _4570_/B _4584_/X vssd1 vssd1 vccd1 vccd1 _4587_/B sky130_fd_sc_hd__a21oi_1
X_7373_ _7373_/A _3662_/Y vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__ebufn_8
XFILLER_89_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6324_ _6324_/A _6327_/A _6324_/C vssd1 vssd1 vccd1 vccd1 _6332_/A sky130_fd_sc_hd__and3_1
X_6255_ _6255_/A _6191_/B vssd1 vssd1 vccd1 vccd1 _6255_/X sky130_fd_sc_hd__or2b_1
X_5206_ hold82/A hold53/A hold87/A vssd1 vssd1 vccd1 vccd1 _5335_/A sky130_fd_sc_hd__and3_1
X_6186_ _6186_/A _6090_/A vssd1 vssd1 vccd1 vccd1 _6186_/X sky130_fd_sc_hd__or2b_1
X_5137_ _5478_/A _5137_/B vssd1 vssd1 vccd1 vccd1 _5289_/B sky130_fd_sc_hd__nand2_1
XFILLER_57_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5068_ _5215_/B _5068_/B vssd1 vssd1 vccd1 vccd1 _5341_/B sky130_fd_sc_hd__and2_1
XFILLER_29_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4019_ _4019_/A _4019_/B vssd1 vssd1 vccd1 vccd1 _4042_/A sky130_fd_sc_hd__xor2_2
XFILLER_44_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold108 hold43/X vssd1 vssd1 vccd1 vccd1 hold108/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold119 _5276_/A vssd1 vssd1 vccd1 vccd1 hold119/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4370_ _4370_/A _4370_/B vssd1 vssd1 vccd1 vccd1 _4370_/Y sky130_fd_sc_hd__nand2_1
XFILLER_98_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _5687_/A _5687_/B _6039_/Y vssd1 vssd1 vccd1 vccd1 _6041_/B sky130_fd_sc_hd__o21a_2
XFILLER_85_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6942_ input6/X _6935_/X _6941_/Y _6939_/X vssd1 vssd1 vccd1 vccd1 _7157_/D sky130_fd_sc_hd__o211a_1
X_6873_ _6873_/A _6873_/B vssd1 vssd1 vccd1 vccd1 _6877_/A sky130_fd_sc_hd__or2_1
X_5824_ _5824_/A vssd1 vssd1 vccd1 vccd1 _6997_/A sky130_fd_sc_hd__buf_2
XFILLER_62_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5755_ _5755_/A _5755_/B vssd1 vssd1 vccd1 vccd1 _5758_/A sky130_fd_sc_hd__nand2_1
X_4706_ _4706_/A _4706_/B vssd1 vssd1 vccd1 vccd1 _4708_/B sky130_fd_sc_hd__nand2_1
X_5686_ _5699_/A _5699_/B vssd1 vssd1 vccd1 vccd1 _5687_/B sky130_fd_sc_hd__nor2_1
X_4637_ _4694_/A vssd1 vssd1 vccd1 vccd1 _7038_/A sky130_fd_sc_hd__clkbuf_2
X_7425_ _7425_/A _3723_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[29] sky130_fd_sc_hd__ebufn_8
X_4568_ _4657_/A _4666_/B vssd1 vssd1 vccd1 vccd1 _4658_/A sky130_fd_sc_hd__nor2_1
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7356_ _7356_/A _3644_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[30] sky130_fd_sc_hd__ebufn_8
X_4499_ _4607_/A vssd1 vssd1 vccd1 vccd1 _4499_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6307_ _6307_/A _6307_/B vssd1 vssd1 vccd1 vccd1 _6307_/Y sky130_fd_sc_hd__nor2_1
X_6238_ _6307_/A _6307_/B vssd1 vssd1 vccd1 vccd1 _6246_/A sky130_fd_sc_hd__xnor2_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ _6169_/A _6169_/B vssd1 vssd1 vccd1 vccd1 _6170_/B sky130_fd_sc_hd__or2_2
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3870_ _5131_/A _7083_/A vssd1 vssd1 vccd1 vccd1 _3978_/A sky130_fd_sc_hd__and2_1
XFILLER_31_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5540_ _5540_/A _5540_/B vssd1 vssd1 vccd1 vccd1 _5543_/A sky130_fd_sc_hd__nand2_1
X_5471_ _5472_/A _5472_/B _5472_/C vssd1 vssd1 vccd1 vccd1 _5531_/B sky130_fd_sc_hd__a21o_1
X_7210_ _7221_/CLK hold92/X vssd1 vssd1 vccd1 vccd1 _7210_/Q sky130_fd_sc_hd__dfxtp_1
X_4422_ _4422_/A _4422_/B vssd1 vssd1 vccd1 vccd1 _4437_/A sky130_fd_sc_hd__xnor2_2
X_7141_ _7151_/CLK hold26/X vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__dfxtp_1
X_4353_ _4353_/A _4353_/B vssd1 vssd1 vccd1 vccd1 _5047_/A sky130_fd_sc_hd__xor2_4
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7072_ _7072_/A _7072_/B vssd1 vssd1 vccd1 vccd1 _7072_/Y sky130_fd_sc_hd__nand2_1
X_4284_ _5347_/A _7183_/Q vssd1 vssd1 vccd1 vccd1 _4285_/B sky130_fd_sc_hd__nor2_1
X_6023_ _6464_/B _6933_/A _6106_/A _6106_/B vssd1 vssd1 vccd1 vccd1 _6023_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_58_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6925_ _7095_/A vssd1 vssd1 vccd1 vccd1 _6954_/B sky130_fd_sc_hd__buf_2
XFILLER_42_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6856_ _6856_/A _6856_/B _6827_/A vssd1 vssd1 vccd1 vccd1 _6856_/X sky130_fd_sc_hd__or3b_1
X_3999_ _7195_/Q _7194_/Q vssd1 vssd1 vccd1 vccd1 _4178_/B sky130_fd_sc_hd__xor2_2
X_6787_ _6751_/A _6753_/Y _6752_/Y vssd1 vssd1 vccd1 vccd1 _6789_/B sky130_fd_sc_hd__a21o_1
X_5807_ _5807_/A _5807_/B vssd1 vssd1 vccd1 vccd1 _5808_/B sky130_fd_sc_hd__nand2_1
XFILLER_50_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5738_ _5787_/A _5737_/C _6589_/A vssd1 vssd1 vccd1 vccd1 _5739_/D sky130_fd_sc_hd__a21o_1
XFILLER_89_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5669_ _5669_/A _5669_/B _5669_/C vssd1 vssd1 vccd1 vccd1 _5673_/A sky130_fd_sc_hd__or3_1
X_7408_ _7408_/A _3703_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[12] sky130_fd_sc_hd__ebufn_8
X_7339_ _7339_/A _3620_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[13] sky130_fd_sc_hd__ebufn_8
X_7304__97 vssd1 vssd1 vccd1 vccd1 _7304__97/HI _7412_/A sky130_fd_sc_hd__conb_1
XFILLER_89_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_95_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4971_ _5146_/B _4971_/B vssd1 vssd1 vccd1 vccd1 _5145_/C sky130_fd_sc_hd__nor2_1
X_3922_ _4011_/A _3922_/B vssd1 vssd1 vccd1 vccd1 _3928_/B sky130_fd_sc_hd__xor2_1
X_6710_ _6710_/A _6611_/A vssd1 vssd1 vccd1 vccd1 _6750_/A sky130_fd_sc_hd__or2b_1
X_3853_ _7211_/Q vssd1 vssd1 vccd1 vccd1 _4003_/A sky130_fd_sc_hd__clkbuf_1
X_6641_ _6640_/A _6641_/B vssd1 vssd1 vccd1 vccd1 _6641_/X sky130_fd_sc_hd__and2b_1
XFILLER_32_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6572_ _6573_/A _6573_/B vssd1 vssd1 vccd1 vccd1 _6596_/B sky130_fd_sc_hd__xor2_1
X_3784_ _3783_/A _3783_/B _3783_/C vssd1 vssd1 vccd1 vccd1 _3785_/C sky130_fd_sc_hd__o21ai_1
X_5523_ _5524_/A _5524_/B vssd1 vssd1 vccd1 vccd1 _5525_/A sky130_fd_sc_hd__nor2_1
X_5454_ _5498_/A _5498_/B vssd1 vssd1 vccd1 vccd1 _5499_/B sky130_fd_sc_hd__xnor2_1
X_4405_ _4405_/A _4405_/B vssd1 vssd1 vccd1 vccd1 _4406_/B sky130_fd_sc_hd__or2_1
X_5385_ _5386_/B _5386_/C _5386_/A vssd1 vssd1 vccd1 vccd1 _5387_/A sky130_fd_sc_hd__o21a_1
X_4336_ _4335_/B _4336_/B vssd1 vssd1 vccd1 vccd1 _4336_/X sky130_fd_sc_hd__and2b_1
X_7124_ _7226_/CLK hold31/X vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__dfxtp_1
XFILLER_101_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7055_ _7055_/A _7072_/B vssd1 vssd1 vccd1 vccd1 _7055_/Y sky130_fd_sc_hd__nand2_1
XFILLER_86_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4267_ _4477_/A _4267_/B vssd1 vssd1 vccd1 vccd1 _4379_/A sky130_fd_sc_hd__nand2_4
X_4198_ _4405_/A _4405_/B vssd1 vssd1 vccd1 vccd1 _4406_/A sky130_fd_sc_hd__nand2_1
XFILLER_86_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6006_ _5935_/Y _5968_/X _5969_/Y _6005_/Y vssd1 vssd1 vccd1 vccd1 _6009_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_55_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6908_ hold30/A _6892_/X _6894_/X hold68/X vssd1 vssd1 vccd1 vccd1 _6908_/X sky130_fd_sc_hd__a22o_1
XFILLER_23_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6839_ _6839_/A _6848_/B vssd1 vssd1 vccd1 vccd1 _6842_/A sky130_fd_sc_hd__xor2_1
XFILLER_23_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5170_ _5804_/A _5168_/X _5169_/Y vssd1 vssd1 vccd1 vccd1 _5171_/C sky130_fd_sc_hd__o21a_1
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4121_ _4025_/A _4025_/B _4120_/X vssd1 vssd1 vccd1 vccd1 _4165_/A sky130_fd_sc_hd__o21ai_2
XFILLER_68_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7295__88 vssd1 vssd1 vccd1 vccd1 _7295__88/HI _7403_/A sky130_fd_sc_hd__conb_1
X_4052_ _7160_/Q _6445_/B vssd1 vssd1 vccd1 vccd1 _4070_/A sky130_fd_sc_hd__and2b_1
Xinput4 io_in[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_2
XFILLER_49_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4954_ _5765_/A _4249_/A _4953_/B vssd1 vssd1 vccd1 vccd1 _4955_/B sky130_fd_sc_hd__a21oi_1
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3905_ _4504_/A _3905_/B vssd1 vssd1 vccd1 vccd1 _3905_/Y sky130_fd_sc_hd__nor2_1
X_4885_ _4889_/A _4889_/B vssd1 vssd1 vccd1 vccd1 _4890_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6624_ _6624_/A _6625_/B vssd1 vssd1 vccd1 vccd1 _6624_/X sky130_fd_sc_hd__or2_1
X_3836_ _7188_/Q vssd1 vssd1 vccd1 vccd1 _6027_/A sky130_fd_sc_hd__buf_2
X_3767_ hold59/X vssd1 vssd1 vccd1 vccd1 _7066_/A sky130_fd_sc_hd__inv_2
X_6555_ _6554_/B _6555_/B vssd1 vssd1 vccd1 vccd1 _6555_/X sky130_fd_sc_hd__and2b_1
X_5506_ _5547_/C _5505_/C _5505_/A vssd1 vssd1 vccd1 vccd1 _5507_/B sky130_fd_sc_hd__a21o_1
X_6486_ _6484_/B _6502_/A _6484_/A vssd1 vssd1 vccd1 vccd1 _6487_/D sky130_fd_sc_hd__a21o_1
X_3698_ _3710_/A vssd1 vssd1 vccd1 vccd1 _3703_/A sky130_fd_sc_hd__buf_8
X_5437_ _5202_/A _5803_/A _6531_/A vssd1 vssd1 vccd1 vccd1 _5438_/A sky130_fd_sc_hd__a21o_1
XFILLER_87_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5368_ _5245_/A _5368_/B vssd1 vssd1 vccd1 vccd1 _5368_/X sky130_fd_sc_hd__and2b_1
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7107_ _3879_/B _7101_/X hold78/X _7099_/X vssd1 vssd1 vccd1 vccd1 hold79/A sky130_fd_sc_hd__o211a_1
X_4319_ _4466_/A _4745_/B _4465_/B vssd1 vssd1 vccd1 vccd1 _4320_/B sky130_fd_sc_hd__a21o_1
X_5299_ _5150_/A _5150_/B _5149_/A vssd1 vssd1 vccd1 vccd1 _5315_/A sky130_fd_sc_hd__a21o_1
XFILLER_101_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7038_ _7038_/A _7038_/B vssd1 vssd1 vccd1 vccd1 _7038_/X sky130_fd_sc_hd__or2_1
XFILLER_74_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4670_ _4670_/A _4670_/B vssd1 vssd1 vccd1 vccd1 _4671_/B sky130_fd_sc_hd__or2_1
X_3621_ _3622_/A vssd1 vssd1 vccd1 vccd1 _3621_/Y sky130_fd_sc_hd__inv_2
X_6340_ _5785_/B _5787_/C _6375_/B vssd1 vssd1 vccd1 vccd1 _6341_/B sky130_fd_sc_hd__mux2_1
XFILLER_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6271_ _6209_/A _6270_/B _6268_/Y vssd1 vssd1 vccd1 vccd1 _6271_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_88_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5222_ _5222_/A _5264_/A vssd1 vssd1 vccd1 vccd1 _5239_/A sky130_fd_sc_hd__xnor2_2
X_5153_ _5154_/A _5154_/B vssd1 vssd1 vccd1 vccd1 _5321_/A sky130_fd_sc_hd__and2_1
XFILLER_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4104_ _6761_/B _4225_/B _6704_/B vssd1 vssd1 vccd1 vccd1 _4372_/B sky130_fd_sc_hd__o21ba_1
XFILLER_96_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5084_ _6034_/A _5085_/B vssd1 vssd1 vccd1 vccd1 _5086_/A sky130_fd_sc_hd__nor2_1
X_4035_ _7223_/Q _6439_/A vssd1 vssd1 vccd1 vccd1 _4036_/C sky130_fd_sc_hd__xnor2_1
XFILLER_64_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5986_ _5986_/A _5986_/B vssd1 vssd1 vccd1 vccd1 _5987_/C sky130_fd_sc_hd__and2_1
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4937_ _4787_/A _4787_/B _4784_/A _4784_/B vssd1 vssd1 vccd1 vccd1 _4940_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_24_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_31 _3739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4868_ _4932_/A _4868_/B vssd1 vssd1 vccd1 vccd1 _4888_/A sky130_fd_sc_hd__nor2_1
XANTENNA_20 _6455_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_42 hold97/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_53 _7045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3819_ hold99/A _3819_/B vssd1 vssd1 vccd1 vccd1 _5145_/A sky130_fd_sc_hd__xnor2_1
XFILLER_20_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6607_ _6415_/B _6607_/B vssd1 vssd1 vccd1 vccd1 _6608_/B sky130_fd_sc_hd__and2b_1
X_4799_ _4799_/A _4799_/B vssd1 vssd1 vccd1 vccd1 _4856_/B sky130_fd_sc_hd__xor2_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6538_ _6538_/A _6538_/B vssd1 vssd1 vccd1 vccd1 _6579_/A sky130_fd_sc_hd__nor2_1
X_6469_ _6475_/D _6473_/A _6472_/B vssd1 vssd1 vccd1 vccd1 _6765_/A sky130_fd_sc_hd__nand3_1
XFILLER_97_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7265__58 vssd1 vssd1 vccd1 vccd1 _7265__58/HI _7364_/A sky130_fd_sc_hd__conb_1
XFILLER_78_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5840_ _5840_/A _5840_/B vssd1 vssd1 vccd1 vccd1 _5841_/A sky130_fd_sc_hd__xnor2_1
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5771_ _5826_/A _5826_/B _5770_/X vssd1 vssd1 vccd1 vccd1 _5774_/B sky130_fd_sc_hd__o21a_1
XFILLER_21_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4722_ _4723_/A _4723_/B vssd1 vssd1 vccd1 vccd1 _4741_/A sky130_fd_sc_hd__nand2_1
XFILLER_21_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4653_ _4653_/A _4653_/B vssd1 vssd1 vccd1 vccd1 _4655_/C sky130_fd_sc_hd__or2_1
X_4584_ _4665_/B _4665_/A vssd1 vssd1 vccd1 vccd1 _4584_/X sky130_fd_sc_hd__and2b_1
X_7372_ _7372_/A _3660_/Y vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__ebufn_8
X_6323_ _6874_/A _6323_/B vssd1 vssd1 vccd1 vccd1 _6353_/A sky130_fd_sc_hd__nand2_1
X_6254_ _6317_/B _6254_/B vssd1 vssd1 vccd1 vccd1 _6258_/A sky130_fd_sc_hd__xnor2_1
X_5205_ hold83/X vssd1 vssd1 vccd1 vccd1 hold82/A sky130_fd_sc_hd__clkbuf_2
X_6185_ _6185_/A _6251_/B vssd1 vssd1 vccd1 vccd1 _6188_/A sky130_fd_sc_hd__xor2_4
XFILLER_84_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5136_ _5478_/A _5137_/B vssd1 vssd1 vccd1 vccd1 _5266_/B sky130_fd_sc_hd__or2_1
X_5067_ _5067_/A _5067_/B _5067_/C vssd1 vssd1 vccd1 vccd1 _5068_/B sky130_fd_sc_hd__nand3_1
X_4018_ _4240_/B _4240_/C _4240_/A vssd1 vssd1 vccd1 vccd1 _4042_/B sky130_fd_sc_hd__a21boi_2
XFILLER_72_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5969_ _5969_/A _5969_/B vssd1 vssd1 vccd1 vccd1 _5969_/Y sky130_fd_sc_hd__nand2_1
XFILLER_40_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold109 _4208_/A vssd1 vssd1 vccd1 vccd1 _7108_/A sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_98_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7314__107 vssd1 vssd1 vccd1 vccd1 _7314__107/HI _7422_/A sky130_fd_sc_hd__conb_1
X_6941_ _6941_/A _6956_/B vssd1 vssd1 vccd1 vccd1 _6941_/Y sky130_fd_sc_hd__nand2_1
X_6872_ _6907_/A vssd1 vssd1 vccd1 vccd1 _6906_/A sky130_fd_sc_hd__clkbuf_2
X_5823_ _5840_/A _5840_/B vssd1 vssd1 vccd1 vccd1 _5823_/X sky130_fd_sc_hd__or2_1
X_5754_ _5773_/A _5754_/B vssd1 vssd1 vccd1 vccd1 _5755_/B sky130_fd_sc_hd__nand2_1
X_4705_ _4760_/A _4760_/B vssd1 vssd1 vccd1 vccd1 _4706_/B sky130_fd_sc_hd__or2b_1
XFILLER_30_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5685_ _5685_/A _5685_/B vssd1 vssd1 vccd1 vccd1 _5699_/B sky130_fd_sc_hd__nor2_2
X_4636_ _4636_/A _4636_/B vssd1 vssd1 vccd1 vccd1 _4717_/A sky130_fd_sc_hd__xnor2_1
X_7424_ _7424_/A _3721_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[28] sky130_fd_sc_hd__ebufn_8
X_7355_ _7355_/A _3643_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[29] sky130_fd_sc_hd__ebufn_8
XFILLER_89_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4567_ _5644_/A _4567_/B vssd1 vssd1 vccd1 vccd1 _4666_/B sky130_fd_sc_hd__nor2_1
X_6306_ _6307_/A _6307_/B vssd1 vssd1 vccd1 vccd1 _6306_/Y sky130_fd_sc_hd__nand2_1
X_4498_ _4498_/A _4498_/B vssd1 vssd1 vccd1 vccd1 _4607_/A sky130_fd_sc_hd__xor2_2
X_6237_ _6170_/A _6170_/B _6236_/X vssd1 vssd1 vccd1 vccd1 _6307_/B sky130_fd_sc_hd__o21ba_1
XFILLER_85_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ _6167_/A _6167_/B _6167_/C vssd1 vssd1 vccd1 vccd1 _6169_/B sky130_fd_sc_hd__a21oi_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5119_ _5119_/A vssd1 vssd1 vccd1 vccd1 _5120_/A sky130_fd_sc_hd__inv_2
XFILLER_57_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6099_ _6192_/A _6192_/B vssd1 vssd1 vccd1 vccd1 _6102_/A sky130_fd_sc_hd__xor2_4
XFILLER_84_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_3_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7151_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_27_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7235__28 vssd1 vssd1 vccd1 vccd1 _7235__28/HI _7334_/A sky130_fd_sc_hd__conb_1
XFILLER_91_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5470_ _5475_/A _5475_/B vssd1 vssd1 vccd1 vccd1 _5472_/C sky130_fd_sc_hd__xnor2_1
X_4421_ _4421_/A _4421_/B vssd1 vssd1 vccd1 vccd1 _4439_/B sky130_fd_sc_hd__xnor2_2
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7140_ _7224_/CLK hold69/X vssd1 vssd1 vccd1 vccd1 hold68/A sky130_fd_sc_hd__dfxtp_1
X_4352_ _5048_/A _4352_/B vssd1 vssd1 vccd1 vccd1 _4353_/B sky130_fd_sc_hd__xnor2_2
XFILLER_98_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7071_ hold99/X _7062_/X _7070_/Y _7060_/X vssd1 vssd1 vccd1 vccd1 _7071_/X sky130_fd_sc_hd__o211a_1
X_4283_ _5812_/A _4325_/B _4282_/X vssd1 vssd1 vccd1 vccd1 _4291_/A sky130_fd_sc_hd__o21ai_2
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6022_ _6022_/A vssd1 vssd1 vccd1 vccd1 _6464_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6924_ hold40/X hold93/X _7117_/B vssd1 vssd1 vccd1 vccd1 _7095_/A sky130_fd_sc_hd__nor3b_1
XFILLER_81_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6855_ _6874_/B _6855_/B vssd1 vssd1 vccd1 vccd1 _6859_/A sky130_fd_sc_hd__and2_1
X_3998_ _7198_/Q _3998_/B vssd1 vssd1 vccd1 vccd1 _4002_/A sky130_fd_sc_hd__xnor2_1
XFILLER_10_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6786_ _6786_/A _6786_/B vssd1 vssd1 vccd1 vccd1 _6789_/A sky130_fd_sc_hd__and2_1
X_5806_ _6523_/A _6160_/A _6061_/B vssd1 vssd1 vccd1 vccd1 _5807_/B sky130_fd_sc_hd__nand3_1
X_5737_ _5737_/A _5787_/A _5737_/C vssd1 vssd1 vccd1 vccd1 _5787_/B sky130_fd_sc_hd__nand3_2
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5668_ _6027_/A _5671_/B _4613_/C vssd1 vssd1 vccd1 vccd1 _5669_/C sky130_fd_sc_hd__a21oi_2
X_7407_ _7407_/A _3702_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[11] sky130_fd_sc_hd__ebufn_8
X_4619_ _4619_/A _4620_/A vssd1 vssd1 vccd1 vccd1 _4692_/B sky130_fd_sc_hd__xnor2_1
X_5599_ _6087_/B _6088_/A vssd1 vssd1 vccd1 vccd1 _5796_/B sky130_fd_sc_hd__nor2_2
X_7338_ _7338_/A _3619_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[12] sky130_fd_sc_hd__ebufn_8
XFILLER_1_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4970_ _5133_/A _5292_/A vssd1 vssd1 vccd1 vccd1 _4971_/B sky130_fd_sc_hd__nor2_1
X_3921_ _3921_/A _3921_/B vssd1 vssd1 vccd1 vccd1 _4008_/A sky130_fd_sc_hd__xor2_1
X_3852_ _3873_/A _3873_/B vssd1 vssd1 vccd1 vccd1 _3877_/C sky130_fd_sc_hd__xor2_2
X_6640_ _6640_/A _6641_/B vssd1 vssd1 vccd1 vccd1 _6650_/B sky130_fd_sc_hd__xnor2_1
XFILLER_32_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6571_ _6571_/A _6571_/B vssd1 vssd1 vccd1 vccd1 _6573_/B sky130_fd_sc_hd__xnor2_1
X_5522_ _5463_/A _5463_/B _5521_/X vssd1 vssd1 vccd1 vccd1 _5524_/B sky130_fd_sc_hd__o21a_1
X_3783_ _3783_/A _3783_/B _3783_/C vssd1 vssd1 vccd1 vccd1 _3785_/B sky130_fd_sc_hd__or3_1
X_5453_ _5352_/A _5352_/B _5351_/A vssd1 vssd1 vccd1 vccd1 _5498_/B sky130_fd_sc_hd__a21bo_1
X_4404_ _4498_/A _4498_/B vssd1 vssd1 vccd1 vccd1 _4407_/B sky130_fd_sc_hd__and2b_1
X_5384_ _5282_/A _5384_/B vssd1 vssd1 vccd1 vccd1 _5386_/C sky130_fd_sc_hd__and2b_1
X_4335_ _4336_/B _4335_/B vssd1 vssd1 vccd1 vccd1 _4445_/B sky130_fd_sc_hd__xnor2_2
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7123_ _7226_/CLK hold49/X vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__dfxtp_1
XFILLER_59_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7054_ hold119/X _6954_/B _7053_/X _7048_/X vssd1 vssd1 vccd1 vccd1 _7198_/D sky130_fd_sc_hd__o211a_1
X_4266_ _5347_/A _7189_/Q vssd1 vssd1 vccd1 vccd1 _4267_/B sky130_fd_sc_hd__or2_2
X_4197_ _4197_/A _4197_/B vssd1 vssd1 vccd1 vccd1 _4405_/B sky130_fd_sc_hd__nor2_1
X_6005_ _6003_/X _6004_/X _5965_/B vssd1 vssd1 vccd1 vccd1 _6005_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_27_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6907_ _6907_/A vssd1 vssd1 vccd1 vccd1 _7116_/A sky130_fd_sc_hd__buf_2
X_6838_ _6812_/A _6812_/B _6837_/Y vssd1 vssd1 vccd1 vccd1 _6848_/B sky130_fd_sc_hd__a21bo_1
XFILLER_23_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6769_ _6769_/A _6797_/B vssd1 vssd1 vccd1 vccd1 _6802_/B sky130_fd_sc_hd__or2_1
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4120_ _4120_/A _4120_/B vssd1 vssd1 vccd1 vccd1 _4120_/X sky130_fd_sc_hd__or2_1
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4051_ _6109_/A _4076_/B vssd1 vssd1 vccd1 vccd1 _4053_/B sky130_fd_sc_hd__nor2_1
Xinput5 io_in[13] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_2
XFILLER_37_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4953_ _5765_/A _4953_/B vssd1 vssd1 vccd1 vccd1 _5127_/A sky130_fd_sc_hd__and2_1
XFILLER_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3904_ _3904_/A vssd1 vssd1 vccd1 vccd1 _4504_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4884_ _4884_/A _4884_/B vssd1 vssd1 vccd1 vccd1 _4889_/B sky130_fd_sc_hd__xor2_1
X_6623_ _6502_/X _6931_/A _6678_/A vssd1 vssd1 vccd1 vccd1 _6625_/B sky130_fd_sc_hd__mux2_1
XFILLER_20_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3835_ _5667_/B vssd1 vssd1 vccd1 vccd1 _4613_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_20_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3766_ _7204_/Q hold70/A vssd1 vssd1 vccd1 vccd1 _4356_/B sky130_fd_sc_hd__xor2_2
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6554_ _6555_/B _6554_/B vssd1 vssd1 vccd1 vccd1 _6579_/B sky130_fd_sc_hd__xnor2_1
X_6485_ _6494_/A _6485_/B vssd1 vssd1 vccd1 vccd1 _6487_/C sky130_fd_sc_hd__or2_1
X_5505_ _5505_/A _5547_/C _5505_/C vssd1 vssd1 vccd1 vccd1 _5507_/A sky130_fd_sc_hd__nand3_1
X_3697_ _3697_/A vssd1 vssd1 vccd1 vccd1 _3697_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5436_ _7175_/Q vssd1 vssd1 vccd1 vccd1 _6531_/A sky130_fd_sc_hd__clkbuf_2
X_5367_ _5367_/A _5367_/B vssd1 vssd1 vccd1 vccd1 _5468_/A sky130_fd_sc_hd__xnor2_1
XFILLER_87_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7106_ hold77/X _7106_/B vssd1 vssd1 vccd1 vccd1 hold78/A sky130_fd_sc_hd__or2_1
X_4318_ hold90/A _5734_/A vssd1 vssd1 vccd1 vccd1 _4465_/B sky130_fd_sc_hd__and2_4
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5298_ _5176_/A _5176_/B _5325_/C vssd1 vssd1 vccd1 vccd1 _5316_/A sky130_fd_sc_hd__o21ai_1
X_4249_ _4249_/A _4506_/B vssd1 vssd1 vccd1 vccd1 _4502_/A sky130_fd_sc_hd__xnor2_1
XFILLER_87_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7037_ _7014_/A _7032_/X _7036_/X _7034_/X vssd1 vssd1 vccd1 vccd1 _7192_/D sky130_fd_sc_hd__o211a_1
XFILLER_19_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3620_ _3622_/A vssd1 vssd1 vccd1 vccd1 _3620_/Y sky130_fd_sc_hd__inv_2
X_6270_ _6270_/A _6270_/B vssd1 vssd1 vccd1 vccd1 _6270_/X sky130_fd_sc_hd__or2_1
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5221_ _5047_/A _5047_/B _5071_/B _5220_/Y vssd1 vssd1 vccd1 vccd1 _5264_/A sky130_fd_sc_hd__a31oi_2
X_5152_ _4995_/A _4995_/B _4979_/A vssd1 vssd1 vccd1 vccd1 _5154_/B sky130_fd_sc_hd__a21o_1
XFILLER_96_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4103_ _5026_/A _4328_/A vssd1 vssd1 vccd1 vccd1 _6704_/B sky130_fd_sc_hd__nor2_2
X_5083_ _5229_/A _5083_/B vssd1 vssd1 vccd1 vccd1 _5085_/B sky130_fd_sc_hd__xnor2_1
X_4034_ _6494_/A vssd1 vssd1 vccd1 vccd1 _6439_/A sky130_fd_sc_hd__buf_2
XFILLER_37_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5985_ _6997_/A _5985_/B vssd1 vssd1 vccd1 vccd1 _5986_/B sky130_fd_sc_hd__or2_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4936_ _4936_/A _4936_/B vssd1 vssd1 vccd1 vccd1 _4940_/A sky130_fd_sc_hd__xnor2_1
XANTENNA_32 _3739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4867_ _4867_/A _4883_/A _4867_/C vssd1 vssd1 vccd1 vccd1 _4868_/B sky130_fd_sc_hd__nor3_1
XANTENNA_10 _7053_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 _6452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_43 hold97/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3818_ _3816_/X _3818_/B vssd1 vssd1 vccd1 vccd1 _3819_/B sky130_fd_sc_hd__and2b_1
X_6606_ _6609_/A _6609_/B vssd1 vssd1 vccd1 vccd1 _6643_/A sky130_fd_sc_hd__xnor2_1
X_4798_ _6931_/A _5937_/B vssd1 vssd1 vccd1 vccd1 _4815_/A sky130_fd_sc_hd__nor2_1
XFILLER_21_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6537_ _6679_/A _6537_/B vssd1 vssd1 vccd1 vccd1 _6538_/B sky130_fd_sc_hd__and2_1
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3749_ _6845_/A vssd1 vssd1 vccd1 vccd1 _5594_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6468_ _6475_/C _6467_/Y _6449_/Y vssd1 vssd1 vccd1 vccd1 _6472_/B sky130_fd_sc_hd__a21o_1
XFILLER_79_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6399_ _6990_/A _6986_/A _6874_/A _6375_/Y vssd1 vssd1 vccd1 vccd1 _6400_/B sky130_fd_sc_hd__o211a_1
X_5419_ _5419_/A _5419_/B vssd1 vssd1 vccd1 vccd1 _5458_/A sky130_fd_sc_hd__nor2_1
XFILLER_101_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5770_ _5770_/A _5770_/B vssd1 vssd1 vccd1 vccd1 _5770_/X sky130_fd_sc_hd__or2_1
X_4721_ _4721_/A vssd1 vssd1 vccd1 vccd1 _6933_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4652_ _4652_/A _4652_/B vssd1 vssd1 vccd1 vccd1 _4653_/B sky130_fd_sc_hd__and2_1
X_4583_ _4580_/A _4580_/B _4671_/A vssd1 vssd1 vccd1 vccd1 _4665_/A sky130_fd_sc_hd__o21ai_2
X_7371_ _7371_/A _3659_/Y vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__ebufn_8
X_6322_ _6369_/B vssd1 vssd1 vccd1 vccd1 _6874_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6253_ _6253_/A _6253_/B vssd1 vssd1 vccd1 vccd1 _6254_/B sky130_fd_sc_hd__nor2_1
XFILLER_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5204_ _5209_/B _5204_/B vssd1 vssd1 vccd1 vccd1 _5213_/A sky130_fd_sc_hd__or2_1
XFILLER_69_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6184_ _6091_/A _6091_/B _6183_/Y vssd1 vssd1 vccd1 vccd1 _6251_/B sky130_fd_sc_hd__a21o_1
X_5135_ _5135_/A _5286_/C vssd1 vssd1 vccd1 vccd1 _5137_/B sky130_fd_sc_hd__xnor2_1
XFILLER_29_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5066_ _5067_/A _5067_/B _5067_/C vssd1 vssd1 vccd1 vccd1 _5215_/B sky130_fd_sc_hd__a21o_1
XFILLER_29_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4017_ _4016_/B _4016_/C _4016_/A vssd1 vssd1 vccd1 vccd1 _4240_/A sky130_fd_sc_hd__a21o_1
XFILLER_84_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5968_ _6007_/A _6007_/B _5967_/Y vssd1 vssd1 vccd1 vccd1 _5968_/X sky130_fd_sc_hd__o21a_1
XFILLER_40_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4919_ _4919_/A _4919_/B vssd1 vssd1 vccd1 vccd1 _4919_/Y sky130_fd_sc_hd__nand2_1
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5899_ _5899_/A _6698_/A vssd1 vssd1 vccd1 vccd1 _5900_/B sky130_fd_sc_hd__and2_1
XFILLER_20_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6940_ input5/X _6935_/X _6938_/Y _6939_/X vssd1 vssd1 vccd1 vccd1 _7156_/D sky130_fd_sc_hd__o211a_1
XFILLER_93_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6871_ _5594_/X hold117/X _5595_/X _6870_/X vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__o211a_1
X_5822_ _5822_/A _5822_/B vssd1 vssd1 vccd1 vccd1 _5845_/B sky130_fd_sc_hd__xnor2_1
XFILLER_34_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5753_ _5773_/A _5754_/B vssd1 vssd1 vccd1 vccd1 _5755_/A sky130_fd_sc_hd__or2_1
X_4704_ _4704_/A _4704_/B vssd1 vssd1 vccd1 vccd1 _4760_/B sky130_fd_sc_hd__xnor2_2
XFILLER_30_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5684_ _5673_/A _5673_/B _5673_/C vssd1 vssd1 vccd1 vccd1 _5685_/B sky130_fd_sc_hd__a21oi_1
X_7423_ _7423_/A _3719_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[27] sky130_fd_sc_hd__ebufn_8
X_4635_ _3802_/Y _4633_/Y _4485_/B _4487_/B _7033_/A vssd1 vssd1 vccd1 vccd1 _4936_/A
+ sky130_fd_sc_hd__a32o_2
X_4566_ _4566_/A _4566_/B vssd1 vssd1 vccd1 vccd1 _4657_/A sky130_fd_sc_hd__or2_1
X_7354_ _7354_/A _3641_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[28] sky130_fd_sc_hd__ebufn_8
X_6305_ _6305_/A _6350_/B vssd1 vssd1 vccd1 vccd1 _6309_/A sky130_fd_sc_hd__xnor2_2
X_4497_ _4497_/A _4497_/B vssd1 vssd1 vccd1 vccd1 _4514_/A sky130_fd_sc_hd__xor2_4
X_6236_ _6156_/A _6236_/B vssd1 vssd1 vccd1 vccd1 _6236_/X sky130_fd_sc_hd__and2b_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6167_ _6167_/A _6167_/B _6167_/C vssd1 vssd1 vccd1 vccd1 _6169_/A sky130_fd_sc_hd__and3_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ _5118_/A _5118_/B vssd1 vssd1 vccd1 vccd1 _5141_/B sky130_fd_sc_hd__nor2_1
XFILLER_84_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6098_ _5893_/A _5893_/B _6097_/Y vssd1 vssd1 vccd1 vccd1 _6192_/B sky130_fd_sc_hd__a21oi_4
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5049_ _3785_/B _5048_/Y _4353_/B _4353_/A vssd1 vssd1 vccd1 vccd1 _5054_/A sky130_fd_sc_hd__a2bb2o_2
XFILLER_25_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4420_ _4407_/X _4496_/B _4495_/A vssd1 vssd1 vccd1 vccd1 _4439_/A sky130_fd_sc_hd__a21o_1
X_4351_ _3783_/B _3783_/C _3783_/A vssd1 vssd1 vccd1 vccd1 _4352_/B sky130_fd_sc_hd__o21ba_1
X_4282_ _5826_/A _6413_/B vssd1 vssd1 vccd1 vccd1 _4282_/X sky130_fd_sc_hd__or2_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7070_ _7070_/A _7072_/B vssd1 vssd1 vccd1 vccd1 _7070_/Y sky130_fd_sc_hd__nand2_1
XFILLER_86_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6021_ _6022_/A _6933_/A _6106_/A vssd1 vssd1 vccd1 vccd1 _6021_/X sky130_fd_sc_hd__and3_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6923_ _6977_/A vssd1 vssd1 vccd1 vccd1 _7116_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6854_ _6854_/A _6854_/B _6854_/C vssd1 vssd1 vccd1 vccd1 _6855_/B sky130_fd_sc_hd__or3_1
XFILLER_35_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3997_ _4022_/A _3997_/B vssd1 vssd1 vccd1 vccd1 _4007_/A sky130_fd_sc_hd__xnor2_1
X_6785_ _6785_/A _6785_/B vssd1 vssd1 vccd1 vccd1 _6786_/B sky130_fd_sc_hd__nand2_1
X_5805_ _6160_/A _5640_/A _6523_/A vssd1 vssd1 vccd1 vccd1 _5807_/A sky130_fd_sc_hd__a21o_1
X_5736_ _5824_/A _5736_/B _5736_/C vssd1 vssd1 vccd1 vccd1 _5736_/X sky130_fd_sc_hd__and3_1
XFILLER_10_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5667_ _7189_/Q _5667_/B vssd1 vssd1 vccd1 vccd1 _5669_/B sky130_fd_sc_hd__and2b_1
X_4618_ _4700_/A _4700_/B _4617_/X vssd1 vssd1 vccd1 vccd1 _4620_/A sky130_fd_sc_hd__o21ba_1
X_7406_ _7406_/A _3701_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[10] sky130_fd_sc_hd__ebufn_8
X_5598_ _5597_/B _5804_/A vssd1 vssd1 vccd1 vccd1 _6088_/A sky130_fd_sc_hd__and2b_1
X_4549_ _4553_/A _4659_/A vssd1 vssd1 vccd1 vccd1 _4550_/B sky130_fd_sc_hd__nand2_1
X_7337_ _7337_/A _3618_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[11] sky130_fd_sc_hd__ebufn_8
XFILLER_89_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6219_ _6219_/A _6219_/B vssd1 vssd1 vccd1 vccd1 _6283_/A sky130_fd_sc_hd__xnor2_2
X_7199_ _7222_/CLK _7199_/D vssd1 vssd1 vccd1 vccd1 _7199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3920_ _3920_/A _3920_/B vssd1 vssd1 vccd1 vccd1 _3931_/A sky130_fd_sc_hd__xnor2_1
XFILLER_17_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3851_ _7196_/Q _3851_/B vssd1 vssd1 vccd1 vccd1 _3873_/B sky130_fd_sc_hd__xnor2_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3782_ _7172_/Q _5736_/B _3781_/X vssd1 vssd1 vccd1 vccd1 _3783_/C sky130_fd_sc_hd__a21boi_1
XFILLER_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6570_ _6978_/A _6592_/B _6569_/A vssd1 vssd1 vccd1 vccd1 _6573_/A sky130_fd_sc_hd__o21a_1
X_5521_ _5521_/A _5521_/B vssd1 vssd1 vccd1 vccd1 _5521_/X sky130_fd_sc_hd__or2_1
X_5452_ _5505_/A _5452_/B vssd1 vssd1 vccd1 vccd1 _5498_/A sky130_fd_sc_hd__nor2_1
X_4403_ _4401_/A _4401_/B _4402_/X vssd1 vssd1 vccd1 vccd1 _4498_/B sky130_fd_sc_hd__o21ai_2
X_5383_ _5383_/A _5383_/B vssd1 vssd1 vccd1 vccd1 _5418_/B sky130_fd_sc_hd__nor2_1
X_4334_ _4334_/A _4334_/B vssd1 vssd1 vccd1 vccd1 _4335_/B sky130_fd_sc_hd__xnor2_1
X_7122_ _7226_/CLK hold20/X vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__dfxtp_1
XFILLER_99_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7053_ _7053_/A _7101_/A vssd1 vssd1 vccd1 vccd1 _7053_/X sky130_fd_sc_hd__or2_1
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6004_ _5971_/X _5998_/Y _6000_/Y _6002_/Y vssd1 vssd1 vccd1 vccd1 _6004_/X sky130_fd_sc_hd__o2bb2a_1
X_4265_ _5098_/A _5098_/B vssd1 vssd1 vccd1 vccd1 _4391_/A sky130_fd_sc_hd__xnor2_2
X_4196_ _4076_/B _4076_/C hold77/A vssd1 vssd1 vccd1 vccd1 _4197_/B sky130_fd_sc_hd__o21a_1
XFILLER_67_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6906_ _6906_/A _6906_/B vssd1 vssd1 vccd1 vccd1 _7147_/D sky130_fd_sc_hd__nor2_1
X_6837_ _6837_/A _6837_/B vssd1 vssd1 vccd1 vccd1 _6837_/Y sky130_fd_sc_hd__nand2_1
X_6768_ _6767_/A _6767_/B _6767_/C vssd1 vssd1 vccd1 vccd1 _6797_/B sky130_fd_sc_hd__a21oi_1
XFILLER_10_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6699_ _6696_/X _6697_/Y _6698_/X vssd1 vssd1 vccd1 vccd1 _6699_/X sky130_fd_sc_hd__a21o_1
X_5719_ _5719_/A _5719_/B vssd1 vssd1 vccd1 vccd1 _5727_/A sky130_fd_sc_hd__xnor2_4
XFILLER_40_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4050_ _6109_/A _4076_/B vssd1 vssd1 vccd1 vccd1 _4054_/A sky130_fd_sc_hd__and2_1
XFILLER_68_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput6 io_in[14] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4952_ _7023_/A _6027_/A vssd1 vssd1 vccd1 vccd1 _4953_/B sky130_fd_sc_hd__and2b_1
XFILLER_51_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4883_ _4883_/A _4883_/B vssd1 vssd1 vccd1 vccd1 _4889_/A sky130_fd_sc_hd__or2_1
X_3903_ _7041_/A _3986_/B _3902_/X vssd1 vssd1 vccd1 vccd1 _3921_/B sky130_fd_sc_hd__a21oi_1
X_6622_ _6622_/A _6622_/B vssd1 vssd1 vccd1 vccd1 _6628_/A sky130_fd_sc_hd__nand2_1
XFILLER_20_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3834_ _4964_/B _3834_/B vssd1 vssd1 vccd1 vccd1 _4950_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3765_ _7201_/Q vssd1 vssd1 vccd1 vccd1 hold70/A sky130_fd_sc_hd__clkbuf_4
X_6553_ _6553_/A _6553_/B vssd1 vssd1 vccd1 vccd1 _6554_/B sky130_fd_sc_hd__xor2_1
X_6484_ _6484_/A _6484_/B _6502_/A vssd1 vssd1 vccd1 vccd1 _6487_/B sky130_fd_sc_hd__nand3_1
X_5504_ _5450_/B _6162_/C _7033_/A vssd1 vssd1 vccd1 vccd1 _5505_/C sky130_fd_sc_hd__o21ai_1
X_3696_ _3697_/A vssd1 vssd1 vccd1 vccd1 _3696_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5435_ _5435_/A _5434_/Y vssd1 vssd1 vccd1 vccd1 _5803_/A sky130_fd_sc_hd__or2b_1
XFILLER_99_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5366_ _5366_/A _5366_/B vssd1 vssd1 vccd1 vccd1 _5367_/B sky130_fd_sc_hd__nor2_1
XFILLER_101_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7105_ hold124/X _7101_/X hold72/X _7099_/X vssd1 vssd1 vccd1 vccd1 hold73/A sky130_fd_sc_hd__o211a_1
XFILLER_59_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5297_ _5382_/A _5382_/B vssd1 vssd1 vccd1 vccd1 _5383_/A sky130_fd_sc_hd__xnor2_1
X_4317_ _4317_/A _4377_/B vssd1 vssd1 vccd1 vccd1 _4321_/A sky130_fd_sc_hd__xnor2_2
X_7286__79 vssd1 vssd1 vccd1 vccd1 _7286__79/HI _7394_/A sky130_fd_sc_hd__conb_1
X_7036_ _7036_/A _7038_/B vssd1 vssd1 vccd1 vccd1 _7036_/X sky130_fd_sc_hd__or2_1
X_4248_ _5722_/A _5667_/B vssd1 vssd1 vccd1 vccd1 _4506_/B sky130_fd_sc_hd__nand2_2
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4179_ _7193_/Q _7192_/Q vssd1 vssd1 vccd1 vccd1 _4531_/B sky130_fd_sc_hd__xor2_4
XFILLER_67_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5220_ _5339_/A _5220_/B vssd1 vssd1 vccd1 vccd1 _5220_/Y sky130_fd_sc_hd__nor2_1
X_5151_ _5151_/A _5151_/B vssd1 vssd1 vccd1 vccd1 _5154_/A sky130_fd_sc_hd__xor2_1
XFILLER_96_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4102_ _4795_/A _4572_/A vssd1 vssd1 vccd1 vccd1 _4328_/A sky130_fd_sc_hd__nand2_4
X_5082_ _4375_/B _4133_/A _5081_/X vssd1 vssd1 vccd1 vccd1 _5083_/B sky130_fd_sc_hd__a21o_1
XFILLER_84_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4033_ _7156_/Q vssd1 vssd1 vccd1 vccd1 _6494_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5984_ _6687_/B vssd1 vssd1 vccd1 vccd1 _6577_/A sky130_fd_sc_hd__clkbuf_2
X_4935_ _4787_/Y _4836_/Y _4838_/X _4839_/Y _4934_/X vssd1 vssd1 vccd1 vccd1 _4935_/X
+ sky130_fd_sc_hd__a2111o_1
X_4866_ _4867_/A _4883_/A _4867_/C vssd1 vssd1 vccd1 vccd1 _4932_/A sky130_fd_sc_hd__o21a_1
XANTENNA_22 _6452_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_11 _6524_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_33 _7099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3817_ _7213_/Q _7199_/Q vssd1 vssd1 vccd1 vccd1 _3818_/B sky130_fd_sc_hd__or2_1
X_4797_ _5991_/A _4796_/X _4328_/A vssd1 vssd1 vccd1 vccd1 _5937_/B sky130_fd_sc_hd__o21ai_4
XANTENNA_44 _6470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6605_ _6605_/A _6605_/B vssd1 vssd1 vccd1 vccd1 _6609_/B sky130_fd_sc_hd__xor2_1
XFILLER_21_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3748_ hold75/X vssd1 vssd1 vccd1 vccd1 _6845_/A sky130_fd_sc_hd__clkbuf_1
X_6536_ _6536_/A _6536_/B vssd1 vssd1 vccd1 vccd1 _6717_/A sky130_fd_sc_hd__xnor2_1
X_6467_ _6480_/A _6821_/A _6588_/A vssd1 vssd1 vccd1 vccd1 _6467_/Y sky130_fd_sc_hd__o21ai_1
X_3679_ _3679_/A vssd1 vssd1 vccd1 vccd1 _3684_/A sky130_fd_sc_hd__buf_6
X_6398_ _6371_/A _6371_/B _6364_/X vssd1 vssd1 vccd1 vccd1 _6400_/A sky130_fd_sc_hd__a21o_1
X_5418_ _5418_/A _5418_/B _5418_/C vssd1 vssd1 vccd1 vccd1 _5419_/B sky130_fd_sc_hd__nor3_1
X_5349_ _5350_/A _5350_/B vssd1 vssd1 vccd1 vccd1 _5351_/A sky130_fd_sc_hd__nand2_1
XFILLER_99_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7019_ _7019_/A _7025_/B vssd1 vssd1 vccd1 vccd1 _7019_/X sky130_fd_sc_hd__or2_1
XFILLER_46_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4720_ _4720_/A _4720_/B vssd1 vssd1 vccd1 vccd1 _4784_/A sky130_fd_sc_hd__xnor2_1
XFILLER_14_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4651_ _4731_/A _4702_/C _4702_/A vssd1 vssd1 vccd1 vccd1 _4703_/A sky130_fd_sc_hd__o21ai_2
X_4582_ _4670_/A _4670_/B vssd1 vssd1 vccd1 vccd1 _4671_/A sky130_fd_sc_hd__nand2_1
X_7370_ _7370_/A _3658_/Y vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__ebufn_8
X_6321_ _6261_/X _6319_/X _6320_/X _6196_/X vssd1 vssd1 vccd1 vccd1 _7132_/D sky130_fd_sc_hd__o211a_1
X_6252_ _6188_/A _6252_/B vssd1 vssd1 vccd1 vccd1 _6253_/B sky130_fd_sc_hd__and2b_1
X_6183_ _6183_/A _6183_/B vssd1 vssd1 vccd1 vccd1 _6183_/Y sky130_fd_sc_hd__nor2_1
X_5203_ _5203_/A _5203_/B vssd1 vssd1 vccd1 vccd1 _5215_/A sky130_fd_sc_hd__nand2_1
XFILLER_69_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5134_ _5287_/B _5134_/B vssd1 vssd1 vccd1 vccd1 _5286_/C sky130_fd_sc_hd__nor2_1
XFILLER_84_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7256__49 vssd1 vssd1 vccd1 vccd1 _7256__49/HI _7355_/A sky130_fd_sc_hd__conb_1
XFILLER_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5065_ _5203_/A _5203_/B vssd1 vssd1 vccd1 vccd1 _5067_/C sky130_fd_sc_hd__xnor2_1
X_4016_ _4016_/A _4016_/B _4016_/C vssd1 vssd1 vccd1 vccd1 _4240_/C sky130_fd_sc_hd__nand3_1
XFILLER_72_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5967_ _5967_/A _5967_/B vssd1 vssd1 vccd1 vccd1 _5967_/Y sky130_fd_sc_hd__nand2_1
X_4918_ _4919_/A _4919_/B vssd1 vssd1 vccd1 vccd1 _4918_/X sky130_fd_sc_hd__or2_1
X_5898_ _5736_/B _5983_/A _5897_/Y vssd1 vssd1 vccd1 vccd1 _5914_/B sky130_fd_sc_hd__o21a_1
X_4849_ hold89/A vssd1 vssd1 vccd1 vccd1 _5913_/A sky130_fd_sc_hd__inv_2
X_6519_ _6487_/X _6566_/A _6512_/X vssd1 vssd1 vccd1 vccd1 _6529_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7270__63 vssd1 vssd1 vccd1 vccd1 _7270__63/HI _7369_/A sky130_fd_sc_hd__conb_1
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6870_ _6877_/B _6869_/X _6261_/A vssd1 vssd1 vccd1 vccd1 _6870_/X sky130_fd_sc_hd__a21o_1
XFILLER_22_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5821_ _5821_/A _5821_/B vssd1 vssd1 vccd1 vccd1 _5822_/B sky130_fd_sc_hd__xor2_1
X_5752_ _5745_/B _5752_/B vssd1 vssd1 vccd1 vccd1 _5754_/B sky130_fd_sc_hd__and2b_1
X_4703_ _4703_/A _4703_/B vssd1 vssd1 vccd1 vccd1 _4760_/A sky130_fd_sc_hd__nand2_1
X_5683_ _5683_/A _5683_/B vssd1 vssd1 vccd1 vccd1 _5699_/A sky130_fd_sc_hd__and2_2
XFILLER_30_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7422_ _7422_/A _3717_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[26] sky130_fd_sc_hd__ebufn_8
X_4634_ _6120_/A vssd1 vssd1 vccd1 vccd1 _7033_/A sky130_fd_sc_hd__buf_2
X_7353_ _7353_/A _3640_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[27] sky130_fd_sc_hd__ebufn_8
X_4565_ _4469_/B _4469_/C _6410_/A vssd1 vssd1 vccd1 vccd1 _4566_/B sky130_fd_sc_hd__a21oi_1
XFILLER_89_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6304_ _6369_/B _6323_/B vssd1 vssd1 vccd1 vccd1 _6350_/B sky130_fd_sc_hd__xor2_1
X_4496_ _4496_/A _4496_/B vssd1 vssd1 vccd1 vccd1 _4604_/A sky130_fd_sc_hd__xnor2_2
X_6235_ _6235_/A _6235_/B vssd1 vssd1 vccd1 vccd1 _6307_/A sky130_fd_sc_hd__xnor2_4
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6166_ _6166_/A _6166_/B vssd1 vssd1 vccd1 vccd1 _6167_/C sky130_fd_sc_hd__xnor2_1
XFILLER_97_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6097_ _6097_/A _6097_/B vssd1 vssd1 vccd1 vccd1 _6097_/Y sky130_fd_sc_hd__nor2_1
X_5117_ _5117_/A _5075_/A vssd1 vssd1 vccd1 vccd1 _5253_/A sky130_fd_sc_hd__or2b_2
X_5048_ _5048_/A vssd1 vssd1 vccd1 vccd1 _5048_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_45_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6999_ _6999_/A _7006_/B vssd1 vssd1 vccd1 vccd1 _6999_/Y sky130_fd_sc_hd__nand2_1
XFILLER_80_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4350_ _4350_/A _5190_/A vssd1 vssd1 vccd1 vccd1 _5048_/A sky130_fd_sc_hd__nor2_2
X_4281_ _5826_/A _6413_/B vssd1 vssd1 vccd1 vccd1 _4325_/B sky130_fd_sc_hd__xnor2_4
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7320__113 vssd1 vssd1 vccd1 vccd1 _7320__113/HI _7428_/A sky130_fd_sc_hd__conb_1
X_6020_ _6020_/A _6020_/B vssd1 vssd1 vccd1 vccd1 _6106_/B sky130_fd_sc_hd__nor2_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6922_ _7052_/A vssd1 vssd1 vccd1 vccd1 _6977_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6853_ _6854_/B _6854_/C _6854_/A vssd1 vssd1 vccd1 vccd1 _6874_/B sky130_fd_sc_hd__o21ai_2
X_5804_ _5804_/A vssd1 vssd1 vccd1 vccd1 _6160_/A sky130_fd_sc_hd__buf_2
XFILLER_50_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3996_ _3996_/A _3996_/B vssd1 vssd1 vccd1 vccd1 _3997_/B sky130_fd_sc_hd__xnor2_1
X_6784_ _6785_/A _6785_/B vssd1 vssd1 vccd1 vccd1 _6786_/A sky130_fd_sc_hd__or2_2
XFILLER_22_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5735_ _5736_/B _5736_/C _5824_/A vssd1 vssd1 vccd1 vccd1 _5745_/A sky130_fd_sc_hd__a21oi_1
X_5666_ _6029_/A vssd1 vssd1 vccd1 vccd1 _5669_/A sky130_fd_sc_hd__inv_2
X_4617_ _4616_/A _4617_/B vssd1 vssd1 vccd1 vccd1 _4617_/X sky130_fd_sc_hd__and2b_1
X_7405_ _7405_/A _3700_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[9] sky130_fd_sc_hd__ebufn_8
X_5597_ _5804_/A _5597_/B vssd1 vssd1 vccd1 vccd1 _6087_/B sky130_fd_sc_hd__and2b_1
X_4548_ _4548_/A _4548_/B vssd1 vssd1 vccd1 vccd1 _4559_/B sky130_fd_sc_hd__xor2_2
X_7336_ _7336_/A _3616_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[10] sky130_fd_sc_hd__ebufn_8
X_4479_ _7202_/Q vssd1 vssd1 vccd1 vccd1 hold91/A sky130_fd_sc_hd__clkbuf_4
XFILLER_89_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6218_ _6216_/Y _6146_/B _6217_/Y vssd1 vssd1 vccd1 vccd1 _6219_/B sky130_fd_sc_hd__a21oi_2
X_7198_ _7221_/CLK _7198_/D vssd1 vssd1 vccd1 vccd1 _7198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6149_ _6149_/A _6149_/B vssd1 vssd1 vccd1 vccd1 _6150_/B sky130_fd_sc_hd__nor2_2
XFILLER_38_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7240__33 vssd1 vssd1 vccd1 vccd1 _7240__33/HI _7339_/A sky130_fd_sc_hd__conb_1
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3850_ _5667_/B _4526_/B vssd1 vssd1 vccd1 vccd1 _3873_/A sky130_fd_sc_hd__nand2_2
XFILLER_32_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3781_ _5619_/B _7168_/Q vssd1 vssd1 vccd1 vccd1 _3781_/X sky130_fd_sc_hd__or2_1
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5520_ _5520_/A _5520_/B vssd1 vssd1 vccd1 vccd1 _5524_/A sky130_fd_sc_hd__xnor2_1
X_5451_ _5228_/B _5483_/C _5348_/S _4285_/A vssd1 vssd1 vccd1 vccd1 _5452_/B sky130_fd_sc_hd__a211oi_1
X_4402_ _7047_/A _4527_/B vssd1 vssd1 vccd1 vccd1 _4402_/X sky130_fd_sc_hd__or2_1
X_5382_ _5382_/A _5382_/B vssd1 vssd1 vccd1 vccd1 _5418_/A sky130_fd_sc_hd__nor2_1
X_4333_ _4436_/A _4435_/B _4332_/Y vssd1 vssd1 vccd1 vccd1 _4336_/B sky130_fd_sc_hd__a21o_1
X_7121_ _7226_/CLK hold22/X vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__dfxtp_1
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4264_ _4491_/A _4491_/B _4263_/X vssd1 vssd1 vccd1 vccd1 _5098_/B sky130_fd_sc_hd__a21oi_2
X_7052_ _7052_/A vssd1 vssd1 vccd1 vccd1 _7101_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6003_ _5971_/X _5998_/Y _6000_/Y _6002_/Y vssd1 vssd1 vccd1 vccd1 _6003_/X sky130_fd_sc_hd__a2bb2o_1
X_4195_ _4195_/A _4195_/B vssd1 vssd1 vccd1 vccd1 _4405_/A sky130_fd_sc_hd__xnor2_1
XFILLER_39_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6905_ hold114/X _6890_/X _6904_/X vssd1 vssd1 vccd1 vccd1 _6906_/B sky130_fd_sc_hd__a21oi_1
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6836_ _6865_/A _6836_/B vssd1 vssd1 vccd1 vccd1 _6839_/A sky130_fd_sc_hd__xor2_1
X_6767_ _6767_/A _6767_/B _6767_/C vssd1 vssd1 vccd1 vccd1 _6769_/A sky130_fd_sc_hd__and3_1
X_5718_ _5718_/A _5718_/B vssd1 vssd1 vccd1 vccd1 _5760_/A sky130_fd_sc_hd__nand2_1
X_3979_ _3979_/A _3979_/B vssd1 vssd1 vccd1 vccd1 _3980_/B sky130_fd_sc_hd__nor2_1
X_6698_ _6698_/A _6698_/B vssd1 vssd1 vccd1 vccd1 _6698_/X sky130_fd_sc_hd__xor2_1
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5649_ _6494_/B _7157_/Q vssd1 vssd1 vccd1 vccd1 _6020_/A sky130_fd_sc_hd__or2b_1
XFILLER_40_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput7 io_in[15] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_2
XFILLER_64_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4951_ _4951_/A _4951_/B vssd1 vssd1 vccd1 vccd1 _4978_/B sky130_fd_sc_hd__nand2_1
X_4882_ _4882_/A _4882_/B vssd1 vssd1 vccd1 vccd1 _4883_/B sky130_fd_sc_hd__and2_1
X_3902_ _4412_/A hold99/A vssd1 vssd1 vccd1 vccd1 _3902_/X sky130_fd_sc_hd__and2_1
X_3833_ _7019_/A _5125_/A _3832_/B vssd1 vssd1 vccd1 vccd1 _3834_/B sky130_fd_sc_hd__o21a_1
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6621_ _6625_/A _6621_/B vssd1 vssd1 vccd1 vccd1 _6622_/B sky130_fd_sc_hd__or2_1
XFILLER_20_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3764_ _3770_/A _3770_/B vssd1 vssd1 vccd1 vccd1 _3801_/A sky130_fd_sc_hd__xnor2_1
X_6552_ _6552_/A _6552_/B vssd1 vssd1 vccd1 vccd1 _6553_/A sky130_fd_sc_hd__nand2_1
XFILLER_20_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6483_ _6483_/A _6483_/B vssd1 vssd1 vccd1 vccd1 _6487_/A sky130_fd_sc_hd__nand2_1
X_3695_ _3697_/A vssd1 vssd1 vccd1 vccd1 _3695_/Y sky130_fd_sc_hd__inv_2
X_5503_ _7033_/A _6209_/A _6162_/C vssd1 vssd1 vccd1 vccd1 _5547_/C sky130_fd_sc_hd__or3_1
X_5434_ _6067_/A _5434_/B vssd1 vssd1 vccd1 vccd1 _5434_/Y sky130_fd_sc_hd__nand2_1
X_7104_ hold71/X _7106_/B vssd1 vssd1 vccd1 vccd1 hold72/A sky130_fd_sc_hd__or2_1
X_5365_ _5241_/B _5365_/B vssd1 vssd1 vccd1 vccd1 _5366_/B sky130_fd_sc_hd__and2b_1
X_4316_ _4316_/A _4316_/B vssd1 vssd1 vccd1 vccd1 _4456_/B sky130_fd_sc_hd__xnor2_1
X_5296_ _5151_/A _5151_/B _5142_/A vssd1 vssd1 vccd1 vccd1 _5382_/B sky130_fd_sc_hd__o21a_1
XFILLER_101_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4247_ _4247_/A _4393_/A vssd1 vssd1 vccd1 vccd1 _4500_/A sky130_fd_sc_hd__xnor2_2
X_7035_ _7011_/A _7032_/X _7033_/X _7034_/X vssd1 vssd1 vccd1 vccd1 _7191_/D sky130_fd_sc_hd__o211a_1
X_4178_ _7197_/Q _4178_/B vssd1 vssd1 vccd1 vccd1 _4182_/A sky130_fd_sc_hd__xnor2_2
XFILLER_55_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_23_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6819_ _5113_/X hold35/X _6817_/Y _6818_/X _3752_/X vssd1 vssd1 vccd1 vccd1 hold36/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_23_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5150_ _5150_/A _5150_/B vssd1 vssd1 vccd1 vccd1 _5151_/B sky130_fd_sc_hd__xnor2_1
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4101_ _5019_/A _4450_/B _6668_/S vssd1 vssd1 vccd1 vccd1 _4225_/B sky130_fd_sc_hd__a21oi_2
X_5081_ _5783_/B _6045_/B _6039_/B vssd1 vssd1 vccd1 vccd1 _5081_/X sky130_fd_sc_hd__and3_1
X_4032_ _7215_/Q _4208_/A vssd1 vssd1 vccd1 vccd1 _4036_/B sky130_fd_sc_hd__or2b_1
XFILLER_56_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5983_ _5983_/A _5983_/B vssd1 vssd1 vccd1 vccd1 _5989_/A sky130_fd_sc_hd__xor2_1
X_4934_ _4934_/A _4934_/B _4934_/C vssd1 vssd1 vccd1 vccd1 _4934_/X sky130_fd_sc_hd__or3_1
X_4865_ _4865_/A _4865_/B vssd1 vssd1 vccd1 vccd1 _4867_/C sky130_fd_sc_hd__and2_1
XANTENNA_23 _6473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_12 _5486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_34 _7099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3816_ _7213_/Q _7199_/Q vssd1 vssd1 vccd1 vccd1 _3816_/X sky130_fd_sc_hd__and2_1
X_4796_ _5596_/A _5596_/B vssd1 vssd1 vccd1 vccd1 _4796_/X sky130_fd_sc_hd__and2_1
X_6604_ _6639_/A _6639_/B _6603_/X vssd1 vssd1 vccd1 vccd1 _6609_/A sky130_fd_sc_hd__a21bo_1
XANTENNA_45 _5091_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3747_ _3747_/A vssd1 vssd1 vccd1 vccd1 _7119_/D sky130_fd_sc_hd__clkbuf_1
X_6535_ _6737_/A _6535_/B vssd1 vssd1 vccd1 vccd1 _6536_/B sky130_fd_sc_hd__xor2_1
XFILLER_21_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6466_ _6466_/A _6466_/B _6821_/A vssd1 vssd1 vccd1 vccd1 _6475_/C sky130_fd_sc_hd__or3_1
X_3678_ _3678_/A vssd1 vssd1 vccd1 vccd1 _3678_/Y sky130_fd_sc_hd__inv_2
X_6397_ _6374_/A _6374_/B _6378_/A _6378_/B vssd1 vssd1 vccd1 vccd1 _6401_/A sky130_fd_sc_hd__o22a_1
X_5417_ _5418_/A _5418_/B _5418_/C vssd1 vssd1 vccd1 vccd1 _5419_/A sky130_fd_sc_hd__o21a_1
XFILLER_99_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5348_ _4289_/A _7053_/A _5348_/S vssd1 vssd1 vccd1 vccd1 _5350_/B sky130_fd_sc_hd__mux2_1
XFILLER_87_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7018_ _7045_/A vssd1 vssd1 vccd1 vccd1 _7018_/X sky130_fd_sc_hd__clkbuf_2
X_5279_ _7055_/A _5280_/B vssd1 vssd1 vccd1 vccd1 _5281_/A sky130_fd_sc_hd__nand2_1
XFILLER_28_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4650_ _4650_/A _4650_/B vssd1 vssd1 vccd1 vccd1 _4702_/A sky130_fd_sc_hd__xor2_1
Xinput10 io_in[18] vssd1 vssd1 vccd1 vccd1 _6891_/B sky130_fd_sc_hd__buf_2
X_4581_ _7001_/A _4914_/B _5871_/A _4468_/A vssd1 vssd1 vccd1 vccd1 _4670_/B sky130_fd_sc_hd__a31o_1
X_6320_ _6391_/A hold10/X vssd1 vssd1 vccd1 vccd1 _6320_/X sky130_fd_sc_hd__or2_1
X_6251_ _6185_/A _6251_/B vssd1 vssd1 vccd1 vccd1 _6253_/A sky130_fd_sc_hd__and2b_1
XFILLER_97_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6182_ _6182_/A _6182_/B vssd1 vssd1 vccd1 vccd1 _6185_/A sky130_fd_sc_hd__xnor2_4
X_5202_ _5202_/A _5330_/A vssd1 vssd1 vccd1 vccd1 _5446_/A sky130_fd_sc_hd__xnor2_4
X_5133_ _5133_/A _7091_/A vssd1 vssd1 vccd1 vccd1 _5134_/B sky130_fd_sc_hd__nor2_1
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5064_ _5209_/B _5064_/B vssd1 vssd1 vccd1 vccd1 _5203_/B sky130_fd_sc_hd__xor2_1
X_4015_ _3844_/X _4821_/B _4016_/B _4245_/A vssd1 vssd1 vccd1 vccd1 _4016_/C sky130_fd_sc_hd__o211ai_1
XFILLER_84_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5966_ _5967_/A _5967_/B vssd1 vssd1 vccd1 vccd1 _6007_/B sky130_fd_sc_hd__nor2_1
XFILLER_13_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4917_ _4899_/Y _4917_/B vssd1 vssd1 vccd1 vccd1 _4919_/A sky130_fd_sc_hd__and2b_1
X_5897_ _6736_/A _5897_/B vssd1 vssd1 vccd1 vccd1 _5897_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4848_ hold90/X vssd1 vssd1 vccd1 vccd1 hold89/A sky130_fd_sc_hd__buf_4
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4779_ _4778_/A _4779_/B vssd1 vssd1 vccd1 vccd1 _4779_/X sky130_fd_sc_hd__and2b_1
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6518_ _6520_/A _6520_/B vssd1 vssd1 vccd1 vccd1 _6529_/A sky130_fd_sc_hd__xnor2_4
X_6449_ _6449_/A _6464_/B vssd1 vssd1 vccd1 vccd1 _6449_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5820_ _5859_/B _5820_/B vssd1 vssd1 vccd1 vccd1 _5865_/A sky130_fd_sc_hd__nor2_1
XFILLER_22_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5751_ _5745_/A _5736_/X _5787_/B _5739_/D vssd1 vssd1 vccd1 vccd1 _5752_/B sky130_fd_sc_hd__a2bb2o_1
X_4702_ _4702_/A _4731_/A _4702_/C vssd1 vssd1 vccd1 vccd1 _4703_/B sky130_fd_sc_hd__or3_1
X_5682_ _5682_/A _5682_/B vssd1 vssd1 vccd1 vccd1 _5683_/B sky130_fd_sc_hd__or2_1
X_7421_ _7421_/A _3714_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[25] sky130_fd_sc_hd__ebufn_8
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4633_ _4633_/A vssd1 vssd1 vccd1 vccd1 _4633_/Y sky130_fd_sc_hd__inv_2
X_4564_ _4564_/A _4564_/B _4564_/C vssd1 vssd1 vccd1 vccd1 _4586_/B sky130_fd_sc_hd__nor3_1
X_7352_ _7352_/A _3639_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[26] sky130_fd_sc_hd__ebufn_8
X_6303_ _6234_/A _6302_/X _6233_/A vssd1 vssd1 vccd1 vccd1 _6323_/B sky130_fd_sc_hd__o21ai_2
X_4495_ _4495_/A _4407_/X vssd1 vssd1 vccd1 vccd1 _4496_/A sky130_fd_sc_hd__or2b_1
X_6234_ _6234_/A _6234_/B vssd1 vssd1 vccd1 vccd1 _6235_/B sky130_fd_sc_hd__xnor2_2
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6165_ _6975_/A _6054_/B _5756_/Y vssd1 vssd1 vccd1 vccd1 _6166_/B sky130_fd_sc_hd__o21a_1
XFILLER_97_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5116_ _5110_/A _5116_/B vssd1 vssd1 vccd1 vccd1 _5257_/A sky130_fd_sc_hd__and2b_1
X_6096_ _6096_/A _6096_/B vssd1 vssd1 vccd1 vccd1 _6192_/A sky130_fd_sc_hd__xnor2_4
X_5047_ _5047_/A _5047_/B vssd1 vssd1 vccd1 vccd1 _5071_/A sky130_fd_sc_hd__nand2_1
XFILLER_27_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6998_ _6679_/A _6993_/X _6997_/X _6995_/X vssd1 vssd1 vccd1 vccd1 _7177_/D sky130_fd_sc_hd__o211a_1
XFILLER_25_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5949_ _6659_/A _5948_/A _5978_/A _5975_/A _5975_/B vssd1 vssd1 vccd1 vccd1 _5955_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_40_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4280_ _5026_/A _4110_/A _4279_/Y vssd1 vssd1 vccd1 vccd1 _6413_/B sky130_fd_sc_hd__o21a_4
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6921_ _6921_/A vssd1 vssd1 vccd1 vccd1 _7052_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6852_ _6852_/A _6852_/B vssd1 vssd1 vccd1 vccd1 _6854_/C sky130_fd_sc_hd__nor2_1
XFILLER_35_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5803_ _5803_/A _5803_/B vssd1 vssd1 vccd1 vccd1 _5815_/B sky130_fd_sc_hd__xnor2_1
X_3995_ _3995_/A _3995_/B vssd1 vssd1 vccd1 vccd1 _3996_/B sky130_fd_sc_hd__nor2_1
X_6783_ _6749_/A _6749_/B _6782_/X vssd1 vssd1 vccd1 vccd1 _6785_/B sky130_fd_sc_hd__a21oi_1
XFILLER_50_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5734_ _5734_/A vssd1 vssd1 vccd1 vccd1 _5824_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5665_ _7186_/Q _7189_/Q vssd1 vssd1 vccd1 vccd1 _6029_/A sky130_fd_sc_hd__or2b_1
X_4616_ _4616_/A _4617_/B vssd1 vssd1 vccd1 vccd1 _4700_/B sky130_fd_sc_hd__xor2_1
X_7404_ _7404_/A _3699_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[8] sky130_fd_sc_hd__ebufn_8
X_7335_ _7335_/A _3615_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[9] sky130_fd_sc_hd__ebufn_8
X_5596_ _5596_/A _5596_/B vssd1 vssd1 vccd1 vccd1 _5602_/A sky130_fd_sc_hd__nand2_2
X_4547_ _4539_/X _4606_/B _4605_/A vssd1 vssd1 vccd1 vccd1 _4559_/A sky130_fd_sc_hd__a21o_1
XFILLER_89_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4478_ _4478_/A _4633_/A vssd1 vssd1 vccd1 vccd1 _4486_/A sky130_fd_sc_hd__or2_1
XFILLER_89_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7197_ _7221_/CLK _7197_/D vssd1 vssd1 vccd1 vccd1 _7197_/Q sky130_fd_sc_hd__dfxtp_2
X_6217_ _6217_/A _6217_/B vssd1 vssd1 vccd1 vccd1 _6217_/Y sky130_fd_sc_hd__nor2_1
X_6148_ _6048_/A _6148_/B vssd1 vssd1 vccd1 vccd1 _6149_/B sky130_fd_sc_hd__and2b_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6079_ _6079_/A _6079_/B vssd1 vssd1 vccd1 vccd1 _6183_/A sky130_fd_sc_hd__xnor2_4
XFILLER_85_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3780_ _5619_/B _7168_/Q vssd1 vssd1 vccd1 vccd1 _5736_/B sky130_fd_sc_hd__nand2_2
XFILLER_12_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5450_ _6162_/C _5450_/B _7053_/A vssd1 vssd1 vccd1 vccd1 _5505_/A sky130_fd_sc_hd__and3b_1
X_4401_ _4401_/A _4401_/B vssd1 vssd1 vccd1 vccd1 _4527_/B sky130_fd_sc_hd__xnor2_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5381_ _5381_/A _5381_/B vssd1 vssd1 vccd1 vccd1 _5528_/A sky130_fd_sc_hd__or2_1
X_4332_ _6421_/A _4332_/B vssd1 vssd1 vccd1 vccd1 _4332_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_3_2_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7226_/CLK
+ sky130_fd_sc_hd__clkbuf_2
X_7120_ _7226_/CLK hold16/X vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__dfxtp_1
X_4263_ _4262_/A _4263_/B vssd1 vssd1 vccd1 vccd1 _4263_/X sky130_fd_sc_hd__and2b_1
X_7051_ _7028_/A _7045_/X _7050_/X _7048_/X vssd1 vssd1 vccd1 vccd1 _7197_/D sky130_fd_sc_hd__o211a_1
XFILLER_59_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6002_ _6002_/A _6002_/B vssd1 vssd1 vccd1 vccd1 _6002_/Y sky130_fd_sc_hd__nand2_1
X_4194_ _4194_/A _4416_/B vssd1 vssd1 vccd1 vccd1 _4195_/B sky130_fd_sc_hd__nor2_1
XFILLER_67_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6904_ hold47/X _6892_/X _6894_/X hold35/X vssd1 vssd1 vccd1 vccd1 _6904_/X sky130_fd_sc_hd__a22o_1
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6835_ _6835_/A _6864_/A vssd1 vssd1 vccd1 vccd1 _6836_/B sky130_fd_sc_hd__xnor2_1
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3978_ _3978_/A _3978_/B _3978_/C vssd1 vssd1 vccd1 vccd1 _3979_/B sky130_fd_sc_hd__nor3_1
X_6766_ _6766_/A _6766_/B vssd1 vssd1 vccd1 vccd1 _6767_/C sky130_fd_sc_hd__xnor2_1
X_5717_ _5717_/A _5872_/A vssd1 vssd1 vccd1 vccd1 _5718_/B sky130_fd_sc_hd__or2_1
XFILLER_10_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6697_ _6690_/A _6693_/Y _6691_/Y vssd1 vssd1 vccd1 vccd1 _6697_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_40_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5648_ _5863_/A _5867_/A _5863_/C vssd1 vssd1 vccd1 vccd1 _5893_/A sky130_fd_sc_hd__a21oi_4
X_5579_ _6264_/A vssd1 vssd1 vccd1 vccd1 _7011_/A sky130_fd_sc_hd__buf_2
XFILLER_65_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7300__93 vssd1 vssd1 vccd1 vccd1 _7300__93/HI _7408_/A sky130_fd_sc_hd__conb_1
XFILLER_58_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput8 io_in[16] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_4
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4950_ _4950_/A _4950_/B vssd1 vssd1 vccd1 vccd1 _4978_/A sky130_fd_sc_hd__nand2_1
XFILLER_51_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4881_ _4884_/A _4884_/B vssd1 vssd1 vccd1 vccd1 _4886_/A sky130_fd_sc_hd__and2b_1
X_3901_ _7210_/Q vssd1 vssd1 vccd1 vccd1 _4412_/A sky130_fd_sc_hd__clkbuf_2
X_3832_ _7019_/A _3832_/B _5125_/A vssd1 vssd1 vccd1 vccd1 _4964_/B sky130_fd_sc_hd__nor3_1
X_6620_ _6620_/A _6620_/B vssd1 vssd1 vccd1 vccd1 _6631_/A sky130_fd_sc_hd__xnor2_2
X_6551_ _6549_/A _6549_/B _6550_/Y vssd1 vssd1 vccd1 vccd1 _6555_/B sky130_fd_sc_hd__a21bo_1
X_3763_ _3785_/A _3763_/B vssd1 vssd1 vccd1 vccd1 _3770_/B sky130_fd_sc_hd__nor2_2
X_5502_ _5444_/A _5444_/B _5442_/A vssd1 vssd1 vccd1 vccd1 _5508_/A sky130_fd_sc_hd__a21oi_1
X_6482_ _6441_/A _6441_/B _6441_/C _6441_/D vssd1 vssd1 vccd1 vccd1 _6491_/B sky130_fd_sc_hd__o22ai_2
X_3694_ _3697_/A vssd1 vssd1 vccd1 vccd1 _3694_/Y sky130_fd_sc_hd__inv_2
X_5433_ _6067_/A _5434_/B vssd1 vssd1 vccd1 vccd1 _5435_/A sky130_fd_sc_hd__nor2_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5364_ _5240_/B _5364_/B vssd1 vssd1 vccd1 vccd1 _5366_/A sky130_fd_sc_hd__and2b_1
X_7103_ _4799_/A _7101_/X _7102_/X _7099_/X vssd1 vssd1 vccd1 vccd1 _7103_/X sky130_fd_sc_hd__o211a_1
X_4315_ _4379_/A _4315_/B vssd1 vssd1 vccd1 vccd1 _4316_/B sky130_fd_sc_hd__xnor2_4
XFILLER_87_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5295_ _5295_/A _5295_/B vssd1 vssd1 vccd1 vccd1 _5382_/A sky130_fd_sc_hd__xnor2_1
X_4246_ _4799_/B _7043_/A vssd1 vssd1 vccd1 vccd1 _4393_/A sky130_fd_sc_hd__nand2_1
X_7034_ _7073_/A vssd1 vssd1 vccd1 vccd1 _7034_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_101_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4177_ _4185_/A _4185_/B vssd1 vssd1 vccd1 vccd1 _4243_/A sky130_fd_sc_hd__xor2_4
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6818_ _6786_/A _6789_/Y _6816_/Y _6879_/A vssd1 vssd1 vccd1 vccd1 _6818_/X sky130_fd_sc_hd__a31o_1
XFILLER_23_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6749_ _6749_/A _6749_/B vssd1 vssd1 vccd1 vccd1 _6750_/C sky130_fd_sc_hd__xnor2_1
XFILLER_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4100_ _4329_/A _4572_/A vssd1 vssd1 vccd1 vccd1 _6668_/S sky130_fd_sc_hd__nor2_1
X_5080_ _5689_/A vssd1 vssd1 vccd1 vccd1 _6034_/A sky130_fd_sc_hd__buf_2
X_4031_ _4039_/A _4039_/B vssd1 vssd1 vccd1 vccd1 _4187_/A sky130_fd_sc_hd__xor2_2
X_7291__84 vssd1 vssd1 vccd1 vccd1 _7291__84/HI _7399_/A sky130_fd_sc_hd__conb_1
X_5982_ _5981_/A _5981_/B _5981_/C vssd1 vssd1 vccd1 vccd1 _5998_/B sky130_fd_sc_hd__a21oi_1
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4933_ _4924_/X _4926_/Y _4932_/Y vssd1 vssd1 vccd1 vccd1 _4934_/C sky130_fd_sc_hd__o21a_1
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4864_ _4864_/A _4864_/B vssd1 vssd1 vccd1 vccd1 _4865_/B sky130_fd_sc_hd__or2_1
XANTENNA_13 _6014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3815_ _3815_/A vssd1 vssd1 vccd1 vccd1 hold99/A sky130_fd_sc_hd__buf_2
XANTENNA_35 _3879_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4795_ _4795_/A _4795_/B vssd1 vssd1 vccd1 vccd1 _5596_/B sky130_fd_sc_hd__or2_1
XANTENNA_46 _6794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_24 _6546_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6603_ _6603_/A _6603_/B _6601_/B vssd1 vssd1 vccd1 vccd1 _6603_/X sky130_fd_sc_hd__or3b_1
X_3746_ _7117_/A _3746_/B vssd1 vssd1 vccd1 vccd1 _3747_/A sky130_fd_sc_hd__and2_1
X_6534_ _6552_/A _6552_/B _6553_/B _6533_/Y vssd1 vssd1 vccd1 vccd1 _6535_/B sky130_fd_sc_hd__a31o_1
X_6465_ _6448_/A _6448_/B _6453_/A vssd1 vssd1 vccd1 vccd1 _6473_/A sky130_fd_sc_hd__o21bai_1
X_3677_ _3678_/A vssd1 vssd1 vccd1 vccd1 _3677_/Y sky130_fd_sc_hd__inv_2
X_5416_ _5416_/A _5416_/B vssd1 vssd1 vccd1 vccd1 _5418_/C sky130_fd_sc_hd__xnor2_1
X_6396_ _6383_/A _6383_/B _6395_/Y vssd1 vssd1 vccd1 vccd1 _6402_/A sky130_fd_sc_hd__a21oi_1
X_5347_ _5347_/A vssd1 vssd1 vccd1 vccd1 _7053_/A sky130_fd_sc_hd__buf_2
XFILLER_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5278_ _5391_/B _5276_/X _5277_/Y _5275_/A vssd1 vssd1 vccd1 vccd1 _5280_/B sky130_fd_sc_hd__a22o_1
XFILLER_101_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7017_ _6997_/A _7005_/X _7016_/X _7007_/X vssd1 vssd1 vccd1 vccd1 _7185_/D sky130_fd_sc_hd__o211a_1
X_4229_ _7179_/Q _7167_/Q vssd1 vssd1 vccd1 vccd1 _4230_/B sky130_fd_sc_hd__or2_1
XFILLER_68_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4580_ _4580_/A _4580_/B vssd1 vssd1 vccd1 vccd1 _4670_/A sky130_fd_sc_hd__xor2_1
Xinput11 io_in[19] vssd1 vssd1 vccd1 vccd1 _6887_/B sky130_fd_sc_hd__clkbuf_4
X_6250_ _6250_/A _6250_/B vssd1 vssd1 vccd1 vccd1 _6317_/B sky130_fd_sc_hd__xor2_1
XFILLER_88_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6181_ _6250_/A _6181_/B vssd1 vssd1 vccd1 vccd1 _6182_/B sky130_fd_sc_hd__and2b_1
X_5201_ _5200_/A _5193_/X _5333_/A _5200_/Y vssd1 vssd1 vccd1 vccd1 _5330_/A sky130_fd_sc_hd__a31o_2
X_5132_ _5133_/A _7091_/A vssd1 vssd1 vccd1 vccd1 _5287_/B sky130_fd_sc_hd__and2_1
XFILLER_96_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5063_ _7072_/A hold58/A _5204_/B vssd1 vssd1 vccd1 vccd1 _5064_/B sky130_fd_sc_hd__o21a_1
X_4014_ _4014_/A _4014_/B vssd1 vssd1 vccd1 vccd1 _4245_/A sky130_fd_sc_hd__xnor2_2
XFILLER_80_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5965_ _5965_/A _5965_/B vssd1 vssd1 vccd1 vccd1 _5967_/B sky130_fd_sc_hd__or2_1
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4916_ _5630_/A _4916_/B vssd1 vssd1 vccd1 vccd1 _5911_/A sky130_fd_sc_hd__nor2_4
X_5896_ _6589_/A vssd1 vssd1 vccd1 vccd1 _6736_/A sky130_fd_sc_hd__buf_2
X_4847_ _4910_/A _4847_/B _4882_/A vssd1 vssd1 vccd1 vccd1 _4902_/A sky130_fd_sc_hd__and3b_1
XFILLER_33_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4778_ _4778_/A _4779_/B vssd1 vssd1 vccd1 vccd1 _4812_/B sky130_fd_sc_hd__xnor2_1
X_6517_ _6724_/A _6724_/B vssd1 vssd1 vccd1 vccd1 _6526_/A sky130_fd_sc_hd__xnor2_4
X_3729_ _3733_/A vssd1 vssd1 vccd1 vccd1 _3729_/Y sky130_fd_sc_hd__inv_2
X_6448_ _6448_/A _6448_/B vssd1 vssd1 vccd1 vccd1 _6452_/A sky130_fd_sc_hd__xnor2_1
X_6379_ _6380_/B _6344_/A vssd1 vssd1 vccd1 vccd1 _6379_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7261__54 vssd1 vssd1 vccd1 vccd1 _7261__54/HI _7360_/A sky130_fd_sc_hd__conb_1
XFILLER_47_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5750_ _6994_/A _5750_/B vssd1 vssd1 vccd1 vccd1 _5773_/A sky130_fd_sc_hd__nor2_1
XFILLER_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4701_ _4704_/B _4704_/A vssd1 vssd1 vccd1 vccd1 _4706_/A sky130_fd_sc_hd__or2b_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5681_ _5689_/A _5681_/B vssd1 vssd1 vccd1 vccd1 _5687_/A sky130_fd_sc_hd__xnor2_2
X_7420_ _7420_/A _3712_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[24] sky130_fd_sc_hd__ebufn_8
X_4632_ _4632_/A _4632_/B vssd1 vssd1 vccd1 vccd1 _4948_/A sky130_fd_sc_hd__xnor2_1
XFILLER_30_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4563_ _4597_/A _4597_/B vssd1 vssd1 vccd1 vccd1 _4600_/A sky130_fd_sc_hd__xnor2_1
X_7351_ _7351_/A _3638_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[25] sky130_fd_sc_hd__ebufn_8
X_4494_ _4494_/A _4494_/B vssd1 vssd1 vccd1 vccd1 _4516_/A sky130_fd_sc_hd__xnor2_4
X_6302_ _6302_/A _6302_/B vssd1 vssd1 vccd1 vccd1 _6302_/X sky130_fd_sc_hd__and2_1
XFILLER_89_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6233_ _6233_/A _6233_/B vssd1 vssd1 vccd1 vccd1 _6234_/B sky130_fd_sc_hd__and2_1
XFILLER_69_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6164_ _6620_/A vssd1 vssd1 vccd1 vccd1 _6975_/A sky130_fd_sc_hd__buf_2
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5115_ _3750_/X hold21/X _3752_/X _5114_/Y vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__o211a_1
X_6095_ _5861_/A _5861_/B _5860_/A vssd1 vssd1 vccd1 vccd1 _6096_/B sky130_fd_sc_hd__a21oi_4
X_5046_ _4165_/A _4165_/B _5045_/X vssd1 vssd1 vccd1 vccd1 _5246_/B sky130_fd_sc_hd__a21bo_1
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6997_ _6997_/A _7011_/B vssd1 vssd1 vccd1 vccd1 _6997_/X sky130_fd_sc_hd__or2_1
XFILLER_53_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5948_ _5948_/A _5948_/B vssd1 vssd1 vccd1 vccd1 _5975_/B sky130_fd_sc_hd__xnor2_1
XFILLER_53_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5879_ _5879_/A _5879_/B vssd1 vssd1 vccd1 vccd1 _5880_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6920_ hold40/A hold93/A _7117_/B vssd1 vssd1 vccd1 vccd1 _6921_/A sky130_fd_sc_hd__or3b_1
XFILLER_62_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6851_ _6990_/A _6851_/B vssd1 vssd1 vccd1 vccd1 _6854_/B sky130_fd_sc_hd__and2_1
X_5802_ _5802_/A _5802_/B vssd1 vssd1 vccd1 vccd1 _5803_/B sky130_fd_sc_hd__nor2_1
X_3994_ _4014_/A _3992_/Y _3993_/Y vssd1 vssd1 vccd1 vccd1 _4022_/A sky130_fd_sc_hd__a21oi_2
X_6782_ _6747_/B _6782_/B vssd1 vssd1 vccd1 vccd1 _6782_/X sky130_fd_sc_hd__and2b_1
XFILLER_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5733_ _6057_/A _6057_/B vssd1 vssd1 vccd1 vccd1 _5748_/A sky130_fd_sc_hd__xnor2_1
X_5664_ _5683_/A _5664_/B vssd1 vssd1 vccd1 vccd1 _6035_/A sky130_fd_sc_hd__xnor2_4
X_7403_ _7403_/A _3697_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[7] sky130_fd_sc_hd__ebufn_8
X_4615_ _4506_/B _4638_/B _4613_/C _4693_/A _4693_/B vssd1 vssd1 vccd1 vccd1 _4617_/B
+ sky130_fd_sc_hd__o32ai_4
X_5595_ _7099_/A vssd1 vssd1 vccd1 vccd1 _5595_/X sky130_fd_sc_hd__clkbuf_2
X_4546_ _4539_/A _4539_/B _4539_/C vssd1 vssd1 vccd1 vccd1 _4605_/A sky130_fd_sc_hd__o21a_1
X_7334_ _7334_/A _3614_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[8] sky130_fd_sc_hd__ebufn_8
X_4477_ _4477_/A _4477_/B vssd1 vssd1 vccd1 vccd1 _4478_/A sky130_fd_sc_hd__and2_1
XFILLER_1_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7196_ _7221_/CLK _7196_/D vssd1 vssd1 vccd1 vccd1 _7196_/Q sky130_fd_sc_hd__dfxtp_2
X_6216_ _6217_/A _6217_/B vssd1 vssd1 vccd1 vccd1 _6216_/Y sky130_fd_sc_hd__nand2_1
XFILLER_58_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6147_ _6041_/B _6147_/B vssd1 vssd1 vccd1 vccd1 _6149_/A sky130_fd_sc_hd__and2b_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6078_ _6078_/A _6078_/B vssd1 vssd1 vccd1 vccd1 _6079_/B sky130_fd_sc_hd__or2_2
X_5029_ _5029_/A _5029_/B vssd1 vssd1 vccd1 vccd1 _5030_/B sky130_fd_sc_hd__xnor2_1
XFILLER_54_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7231__24 vssd1 vssd1 vccd1 vccd1 _7231__24/HI _7330_/A sky130_fd_sc_hd__conb_1
XFILLER_32_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4400_ _4400_/A vssd1 vssd1 vccd1 vccd1 _7047_/A sky130_fd_sc_hd__inv_2
X_5380_ _5380_/A _5380_/B vssd1 vssd1 vccd1 vccd1 _5472_/A sky130_fd_sc_hd__or2_1
XFILLER_99_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4331_ _6421_/A _4332_/B vssd1 vssd1 vccd1 vccd1 _4435_/B sky130_fd_sc_hd__nand2_1
X_4262_ _4262_/A _4263_/B vssd1 vssd1 vccd1 vccd1 _4491_/B sky130_fd_sc_hd__xnor2_4
X_7050_ hold99/X _7059_/B vssd1 vssd1 vccd1 vccd1 _7050_/X sky130_fd_sc_hd__or2_1
XFILLER_101_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6001_ _6001_/A _6001_/B vssd1 vssd1 vccd1 vccd1 _6002_/B sky130_fd_sc_hd__or2_1
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4193_ _5131_/A _4193_/B vssd1 vssd1 vccd1 vccd1 _4416_/B sky130_fd_sc_hd__xnor2_2
XFILLER_39_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6903_ _6906_/A _6903_/B vssd1 vssd1 vccd1 vccd1 _7146_/D sky130_fd_sc_hd__nor2_1
XFILLER_62_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6834_ _6808_/A _6808_/B _6833_/X vssd1 vssd1 vccd1 vccd1 _6864_/A sky130_fd_sc_hd__a21oi_1
X_6765_ _6765_/A _6765_/B vssd1 vssd1 vccd1 vccd1 _6766_/B sky130_fd_sc_hd__nand2_1
X_3977_ _3978_/B _3978_/C _3978_/A vssd1 vssd1 vccd1 vccd1 _3979_/A sky130_fd_sc_hd__o21a_1
X_5716_ _5716_/A _5716_/B vssd1 vssd1 vccd1 vccd1 _5731_/B sky130_fd_sc_hd__xnor2_2
X_6696_ _6691_/A _6691_/B _6691_/Y _6692_/X _6695_/X vssd1 vssd1 vccd1 vccd1 _6696_/X
+ sky130_fd_sc_hd__o2111a_1
X_5647_ _5647_/A _5647_/B vssd1 vssd1 vccd1 vccd1 _5863_/C sky130_fd_sc_hd__xor2_2
X_5578_ _5559_/A _5578_/B vssd1 vssd1 vccd1 vccd1 _5578_/X sky130_fd_sc_hd__and2b_1
X_4529_ _4611_/A _4529_/B vssd1 vssd1 vccd1 vccd1 _4608_/A sky130_fd_sc_hd__xnor2_1
XFILLER_49_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7297__90 vssd1 vssd1 vccd1 vccd1 _7297__90/HI _7405_/A sky130_fd_sc_hd__conb_1
X_7179_ _7183_/CLK _7179_/D vssd1 vssd1 vccd1 vccd1 _7179_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7310__103 vssd1 vssd1 vccd1 vccd1 _7310__103/HI _7418_/A sky130_fd_sc_hd__conb_1
XFILLER_41_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput9 io_in[17] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_2
XFILLER_91_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4880_ _4876_/A _4895_/B _4892_/A vssd1 vssd1 vccd1 vccd1 _4884_/B sky130_fd_sc_hd__o21ai_2
X_3900_ _7210_/Q _7197_/Q vssd1 vssd1 vccd1 vccd1 _3986_/B sky130_fd_sc_hd__xor2_2
XFILLER_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3831_ _7188_/Q _5674_/B vssd1 vssd1 vccd1 vccd1 _5125_/A sky130_fd_sc_hd__nand2_2
X_3762_ _3761_/C _3761_/B _3805_/A vssd1 vssd1 vccd1 vccd1 _3763_/B sky130_fd_sc_hd__a21boi_1
X_6550_ _6575_/A _6575_/B vssd1 vssd1 vccd1 vccd1 _6550_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5501_ _5415_/A _5501_/B vssd1 vssd1 vccd1 vccd1 _5510_/B sky130_fd_sc_hd__and2b_1
X_6481_ _6481_/A _6481_/B vssd1 vssd1 vccd1 vccd1 _6514_/A sky130_fd_sc_hd__xor2_2
X_3693_ _3697_/A vssd1 vssd1 vccd1 vccd1 _3693_/Y sky130_fd_sc_hd__inv_2
X_5432_ _5432_/A _5782_/B vssd1 vssd1 vccd1 vccd1 _5434_/B sky130_fd_sc_hd__nand2_1
XFILLER_99_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5363_ _5464_/A _5464_/B vssd1 vssd1 vccd1 vccd1 _5367_/A sky130_fd_sc_hd__xnor2_1
X_7102_ _7102_/A _7106_/B vssd1 vssd1 vccd1 vccd1 _7102_/X sky130_fd_sc_hd__or2_1
X_4314_ _4469_/B _4452_/B _4313_/Y vssd1 vssd1 vccd1 vccd1 _4316_/A sky130_fd_sc_hd__o21a_1
XFILLER_101_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5294_ _5294_/A _5294_/B vssd1 vssd1 vccd1 vccd1 _5295_/B sky130_fd_sc_hd__xnor2_1
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4245_ _4245_/A _4245_/B vssd1 vssd1 vccd1 vccd1 _4257_/A sky130_fd_sc_hd__xnor2_2
X_7033_ _7033_/A _7038_/B vssd1 vssd1 vccd1 vccd1 _7033_/X sky130_fd_sc_hd__or2_1
X_4176_ _4176_/A _4176_/B vssd1 vssd1 vccd1 vccd1 _4185_/B sky130_fd_sc_hd__xnor2_2
XFILLER_55_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6817_ _6786_/A _6789_/Y _6816_/Y vssd1 vssd1 vccd1 vccd1 _6817_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6748_ _6828_/A _6584_/B _6413_/B vssd1 vssd1 vccd1 vccd1 _6749_/B sky130_fd_sc_hd__o21ba_1
XFILLER_51_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6679_ _6679_/A _6679_/B vssd1 vssd1 vccd1 vccd1 _6688_/A sky130_fd_sc_hd__xnor2_1
XFILLER_76_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4030_ _4189_/A _4189_/B vssd1 vssd1 vccd1 vccd1 _4039_/B sky130_fd_sc_hd__nor2_1
XFILLER_37_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5981_ _5981_/A _5981_/B _5981_/C vssd1 vssd1 vccd1 vccd1 _6000_/B sky130_fd_sc_hd__and3_1
X_4932_ _4932_/A _4932_/B vssd1 vssd1 vccd1 vccd1 _4932_/Y sky130_fd_sc_hd__nor2_1
X_4863_ _4882_/A _4882_/B vssd1 vssd1 vccd1 vccd1 _4883_/A sky130_fd_sc_hd__nor2_1
XANTENNA_14 _6029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6602_ _6603_/B _6602_/B vssd1 vssd1 vccd1 vccd1 _6639_/B sky130_fd_sc_hd__xnor2_2
XANTENNA_36 _3879_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3814_ _5765_/A vssd1 vssd1 vccd1 vccd1 _7019_/A sky130_fd_sc_hd__clkbuf_4
X_4794_ _4794_/A _4795_/B vssd1 vssd1 vccd1 vccd1 _5596_/A sky130_fd_sc_hd__nand2_1
XANTENNA_47 _7114_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_25 _6802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3745_ _7020_/A vssd1 vssd1 vccd1 vccd1 _7117_/A sky130_fd_sc_hd__clkbuf_4
X_6533_ _6540_/A _6533_/B vssd1 vssd1 vccd1 vccd1 _6533_/Y sky130_fd_sc_hd__nor2_1
X_6464_ _6464_/A _6464_/B _6496_/B vssd1 vssd1 vccd1 vccd1 _6475_/D sky130_fd_sc_hd__or3_1
X_3676_ _3678_/A vssd1 vssd1 vccd1 vccd1 _3676_/Y sky130_fd_sc_hd__inv_2
X_5415_ _5415_/A _5501_/B vssd1 vssd1 vccd1 vccd1 _5416_/B sky130_fd_sc_hd__xnor2_1
X_6395_ _6395_/A _6395_/B vssd1 vssd1 vccd1 vccd1 _6395_/Y sky130_fd_sc_hd__nor2_1
X_5346_ _5161_/A _5166_/B _5483_/C vssd1 vssd1 vccd1 vccd1 _5350_/A sky130_fd_sc_hd__o21ai_1
XFILLER_87_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5277_ _5391_/B _5277_/B vssd1 vssd1 vccd1 vccd1 _5277_/Y sky130_fd_sc_hd__nor2_1
XFILLER_87_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7016_ _7016_/A _7025_/B vssd1 vssd1 vccd1 vccd1 _7016_/X sky130_fd_sc_hd__or2_1
X_4228_ _4317_/A hold90/A vssd1 vssd1 vccd1 vccd1 _5750_/B sky130_fd_sc_hd__nand2_8
X_7267__60 vssd1 vssd1 vccd1 vccd1 _7267__60/HI _7366_/A sky130_fd_sc_hd__conb_1
X_4159_ _4159_/A _4159_/B vssd1 vssd1 vccd1 vccd1 _4162_/A sky130_fd_sc_hd__xor2_1
XFILLER_28_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput12 io_in[20] vssd1 vssd1 vccd1 vccd1 _6887_/A sky130_fd_sc_hd__clkbuf_2
X_6180_ _6180_/A _6180_/B _6180_/C vssd1 vssd1 vccd1 vccd1 _6181_/B sky130_fd_sc_hd__or3_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5200_ _5200_/A _5430_/A vssd1 vssd1 vccd1 vccd1 _5200_/Y sky130_fd_sc_hd__nor2_1
XFILLER_96_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5131_ _5131_/A vssd1 vssd1 vccd1 vccd1 _7091_/A sky130_fd_sc_hd__buf_2
XFILLER_57_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5062_ _7070_/A _7202_/Q _5062_/C vssd1 vssd1 vccd1 vccd1 _5204_/B sky130_fd_sc_hd__or3_1
XFILLER_96_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4013_ _4506_/C vssd1 vssd1 vccd1 vccd1 _4821_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_84_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5964_ _5969_/A _5969_/B vssd1 vssd1 vccd1 vccd1 _5965_/B sky130_fd_sc_hd__nor2_1
X_4915_ _5734_/A _5880_/B vssd1 vssd1 vccd1 vccd1 _4916_/B sky130_fd_sc_hd__nor2_1
X_5895_ _5895_/A _5897_/B vssd1 vssd1 vccd1 vccd1 _5914_/A sky130_fd_sc_hd__xor2_1
XFILLER_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4846_ _5829_/B _6409_/B vssd1 vssd1 vccd1 vccd1 _4882_/A sky130_fd_sc_hd__nand2_1
X_4777_ _4814_/A _4814_/B _4776_/X vssd1 vssd1 vccd1 vccd1 _4779_/B sky130_fd_sc_hd__a21bo_1
X_6516_ _6797_/A _6566_/A _6490_/X _6515_/X vssd1 vssd1 vccd1 vccd1 _6724_/B sky130_fd_sc_hd__a211oi_4
X_3728_ _3734_/A vssd1 vssd1 vccd1 vccd1 _3733_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6447_ _6679_/B _6434_/B _6507_/B vssd1 vssd1 vccd1 vccd1 _6448_/B sky130_fd_sc_hd__a21oi_1
X_3659_ _3660_/A vssd1 vssd1 vccd1 vccd1 _3659_/Y sky130_fd_sc_hd__inv_2
X_6378_ _6378_/A _6378_/B vssd1 vssd1 vccd1 vccd1 _6395_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5329_ _5784_/A vssd1 vssd1 vccd1 vccd1 _6539_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_57_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4700_ _4700_/A _4700_/B vssd1 vssd1 vccd1 vccd1 _4704_/A sky130_fd_sc_hd__xor2_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5680_ _6035_/A _6035_/B vssd1 vssd1 vccd1 vccd1 _5681_/B sky130_fd_sc_hd__xor2_2
X_4631_ _5108_/A _5108_/B vssd1 vssd1 vccd1 vccd1 _4632_/B sky130_fd_sc_hd__xor2_1
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4562_ _4562_/A _4562_/B vssd1 vssd1 vccd1 vccd1 _4597_/B sky130_fd_sc_hd__xor2_1
X_7350_ _7350_/A _3637_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[24] sky130_fd_sc_hd__ebufn_8
X_4493_ _4493_/A _4493_/B vssd1 vssd1 vccd1 vccd1 _4601_/A sky130_fd_sc_hd__nor2_1
X_6301_ _6301_/A vssd1 vssd1 vccd1 vccd1 _6369_/B sky130_fd_sc_hd__clkbuf_2
X_6232_ _6302_/A _6302_/B vssd1 vssd1 vccd1 vccd1 _6233_/B sky130_fd_sc_hd__nand2_1
XFILLER_97_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6163_ _6234_/A _6163_/B vssd1 vssd1 vccd1 vccd1 _6166_/A sky130_fd_sc_hd__and2_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5114_ _5111_/X _5257_/B _5113_/X vssd1 vssd1 vccd1 vccd1 _5114_/Y sky130_fd_sc_hd__o21ai_1
X_6094_ _6189_/A _6189_/B vssd1 vssd1 vccd1 vccd1 _6096_/A sky130_fd_sc_hd__xnor2_4
XFILLER_84_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5045_ _5045_/A _4166_/A vssd1 vssd1 vccd1 vccd1 _5045_/X sky130_fd_sc_hd__or2b_1
X_7237__30 vssd1 vssd1 vccd1 vccd1 _7237__30/HI _7336_/A sky130_fd_sc_hd__conb_1
XFILLER_38_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6996_ _6971_/A _6993_/X _6994_/Y _6995_/X vssd1 vssd1 vccd1 vccd1 _7176_/D sky130_fd_sc_hd__o211a_1
XFILLER_53_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5947_ _6659_/A _5978_/A _5945_/A vssd1 vssd1 vccd1 vccd1 _5948_/B sky130_fd_sc_hd__o21ba_1
XFILLER_13_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5878_ _5879_/B vssd1 vssd1 vccd1 vccd1 _5878_/Y sky130_fd_sc_hd__inv_2
X_4829_ _4830_/A _4830_/B vssd1 vssd1 vccd1 vccd1 _4927_/B sky130_fd_sc_hd__and2_1
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6850_ _6850_/A _6850_/B vssd1 vssd1 vccd1 vccd1 _6862_/B sky130_fd_sc_hd__nor2_1
XFILLER_35_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6781_ _6793_/A _6793_/B vssd1 vssd1 vccd1 vccd1 _6785_/A sky130_fd_sc_hd__xnor2_1
XFILLER_35_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5801_ _5801_/A _5801_/B vssd1 vssd1 vccd1 vccd1 _5802_/B sky130_fd_sc_hd__nor2_1
XFILLER_50_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3993_ _4504_/A _3993_/B vssd1 vssd1 vccd1 vccd1 _3993_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5732_ _5759_/A _5759_/B _5731_/X vssd1 vssd1 vccd1 vccd1 _6057_/B sky130_fd_sc_hd__a21oi_2
X_5663_ _6020_/B _5663_/B vssd1 vssd1 vccd1 vccd1 _5664_/B sky130_fd_sc_hd__xor2_4
X_4614_ _7023_/A _4503_/Y _4614_/S vssd1 vssd1 vccd1 vccd1 _4693_/B sky130_fd_sc_hd__mux2_2
X_5594_ _5594_/A vssd1 vssd1 vccd1 vccd1 _5594_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7402_ _7402_/A _3696_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[6] sky130_fd_sc_hd__ebufn_8
X_4545_ _4545_/A vssd1 vssd1 vccd1 vccd1 _4606_/B sky130_fd_sc_hd__inv_2
X_7333_ _7333_/A _3613_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[7] sky130_fd_sc_hd__ebufn_8
X_4476_ _7191_/Q vssd1 vssd1 vccd1 vccd1 _6120_/A sky130_fd_sc_hd__buf_2
X_7195_ _7221_/CLK _7195_/D vssd1 vssd1 vccd1 vccd1 _7195_/Q sky130_fd_sc_hd__dfxtp_1
X_6215_ _6215_/A _6215_/B vssd1 vssd1 vccd1 vccd1 _6219_/A sky130_fd_sc_hd__xnor2_2
XFILLER_85_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6146_ _6146_/A _6146_/B vssd1 vssd1 vccd1 vccd1 _6223_/B sky130_fd_sc_hd__xnor2_4
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6077_ _6076_/A _6076_/B _6076_/C vssd1 vssd1 vccd1 vccd1 _6078_/B sky130_fd_sc_hd__o21a_1
X_5028_ _5171_/B _5028_/B vssd1 vssd1 vccd1 vccd1 _5029_/B sky130_fd_sc_hd__and2_1
XFILLER_26_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6979_ _7007_/A vssd1 vssd1 vccd1 vccd1 _6979_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4330_ _4330_/A _5854_/A vssd1 vssd1 vccd1 vccd1 _4332_/B sky130_fd_sc_hd__or2_1
XFILLER_99_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4261_ _4494_/A _4494_/B _4260_/X vssd1 vssd1 vccd1 vccd1 _4263_/B sky130_fd_sc_hd__a21bo_2
X_6000_ _6000_/A _6000_/B vssd1 vssd1 vccd1 vccd1 _6000_/Y sky130_fd_sc_hd__nor2_1
X_4192_ _3879_/B _4726_/B _4540_/B vssd1 vssd1 vccd1 vccd1 _4194_/A sky130_fd_sc_hd__a21oi_1
XFILLER_79_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6902_ hold37/X _6890_/X _6901_/X vssd1 vssd1 vccd1 vccd1 _6903_/B sky130_fd_sc_hd__a21oi_1
XFILLER_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6833_ _6807_/B _6833_/B vssd1 vssd1 vccd1 vccd1 _6833_/X sky130_fd_sc_hd__and2b_1
XFILLER_62_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3976_ _3943_/B _4026_/A vssd1 vssd1 vccd1 vccd1 _3978_/C sky130_fd_sc_hd__and2b_1
X_6764_ _6978_/A _6736_/B _6763_/Y vssd1 vssd1 vccd1 vccd1 _6772_/A sky130_fd_sc_hd__a21o_1
X_6695_ _6950_/A _6693_/Y _6694_/X _6688_/B vssd1 vssd1 vccd1 vccd1 _6695_/X sky130_fd_sc_hd__a211o_1
X_5715_ _5715_/A _5715_/B vssd1 vssd1 vccd1 vccd1 _5716_/A sky130_fd_sc_hd__nand2_1
X_5646_ _5936_/A _6691_/A _4744_/B vssd1 vssd1 vccd1 vccd1 _5647_/B sky130_fd_sc_hd__a21o_2
X_5577_ _5575_/A _5575_/B _5564_/A vssd1 vssd1 vccd1 vccd1 _5589_/A sky130_fd_sc_hd__o21ai_1
X_4528_ _4611_/A _4529_/B vssd1 vssd1 vccd1 vccd1 _4539_/A sky130_fd_sc_hd__and2_1
XFILLER_2_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4459_ _7176_/Q _5167_/A vssd1 vssd1 vccd1 vccd1 _4469_/C sky130_fd_sc_hd__or2_1
XFILLER_58_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7178_ _7225_/CLK _7178_/D vssd1 vssd1 vccd1 vccd1 _7178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6129_ _6129_/A _6129_/B vssd1 vssd1 vccd1 vccd1 _6129_/Y sky130_fd_sc_hd__nand2_1
XFILLER_65_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3830_ _7187_/Q vssd1 vssd1 vccd1 vccd1 _5674_/B sky130_fd_sc_hd__buf_2
XFILLER_32_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3761_ _3805_/A _3761_/B _3761_/C vssd1 vssd1 vccd1 vccd1 _3785_/A sky130_fd_sc_hd__and3b_1
X_5500_ _5414_/B _5500_/B vssd1 vssd1 vccd1 vccd1 _5510_/A sky130_fd_sc_hd__and2b_1
X_6480_ _6480_/A _6480_/B _6480_/C vssd1 vssd1 vccd1 vccd1 _6566_/A sky130_fd_sc_hd__and3_2
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3692_ _3710_/A vssd1 vssd1 vccd1 vccd1 _3697_/A sky130_fd_sc_hd__buf_12
XFILLER_9_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5431_ _5784_/A _6575_/A vssd1 vssd1 vccd1 vccd1 _5782_/B sky130_fd_sc_hd__nand2_1
X_5362_ _5242_/A _5242_/B _5361_/Y vssd1 vssd1 vccd1 vccd1 _5464_/B sky130_fd_sc_hd__o21a_1
XFILLER_99_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4313_ _4460_/A _5871_/A vssd1 vssd1 vccd1 vccd1 _4313_/Y sky130_fd_sc_hd__nand2_1
X_7101_ _7101_/A vssd1 vssd1 vccd1 vccd1 _7101_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_99_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7032_ _7045_/A vssd1 vssd1 vccd1 vccd1 _7032_/X sky130_fd_sc_hd__clkbuf_2
X_5293_ _5391_/A _5293_/B vssd1 vssd1 vccd1 vccd1 _5294_/B sky130_fd_sc_hd__nand2_1
XFILLER_101_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4244_ _3844_/X _4821_/B _4016_/B vssd1 vssd1 vccd1 vccd1 _4245_/B sky130_fd_sc_hd__o21a_1
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4175_ _4857_/B _7043_/A _4247_/A _4174_/X vssd1 vssd1 vccd1 vccd1 _4185_/A sky130_fd_sc_hd__a31o_2
XFILLER_67_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6816_ _6840_/A _6816_/B vssd1 vssd1 vccd1 vccd1 _6816_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6747_ _6782_/B _6747_/B vssd1 vssd1 vccd1 vccd1 _6749_/A sky130_fd_sc_hd__xnor2_1
X_3959_ _5016_/A _6941_/A vssd1 vssd1 vccd1 vccd1 _3960_/D sky130_fd_sc_hd__or2_1
X_6678_ _6678_/A vssd1 vssd1 vccd1 vccd1 _6926_/A sky130_fd_sc_hd__clkbuf_2
X_5629_ _5623_/Y _5897_/B _5628_/Y vssd1 vssd1 vccd1 vccd1 _5869_/B sky130_fd_sc_hd__a21oi_2
XFILLER_78_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5980_ _5999_/B _5980_/B vssd1 vssd1 vccd1 vccd1 _5981_/C sky130_fd_sc_hd__xnor2_1
X_4931_ _4931_/A _4931_/B vssd1 vssd1 vccd1 vccd1 _4934_/B sky130_fd_sc_hd__nor2_1
XFILLER_64_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4862_ _4867_/A _4862_/B vssd1 vssd1 vccd1 vccd1 _4882_/B sky130_fd_sc_hd__or2_1
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3813_ _5667_/B vssd1 vssd1 vccd1 vccd1 _5765_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_60_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6601_ _6603_/A _6601_/B vssd1 vssd1 vccd1 vccd1 _6602_/B sky130_fd_sc_hd__and2b_1
X_4793_ _6507_/A vssd1 vssd1 vccd1 vccd1 _6931_/A sky130_fd_sc_hd__buf_2
XANTENNA_48 _7059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_37 _4553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_26 _6889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_15 _5699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6532_ _6540_/A _6533_/B vssd1 vssd1 vccd1 vccd1 _6553_/B sky130_fd_sc_hd__xor2_1
X_3744_ _7020_/A vssd1 vssd1 vccd1 vccd1 _7226_/D sky130_fd_sc_hd__clkbuf_2
X_6463_ _6485_/B _6494_/B vssd1 vssd1 vccd1 vccd1 _6496_/B sky130_fd_sc_hd__xnor2_2
X_3675_ _3678_/A vssd1 vssd1 vccd1 vccd1 _3675_/Y sky130_fd_sc_hd__inv_2
X_5414_ _5500_/B _5414_/B vssd1 vssd1 vccd1 vccd1 _5501_/B sky130_fd_sc_hd__xnor2_1
X_6394_ _6390_/A _6390_/B _6393_/X vssd1 vssd1 vccd1 vccd1 _6403_/A sky130_fd_sc_hd__a21o_1
X_5345_ _5450_/B _5232_/B _5231_/B vssd1 vssd1 vccd1 vccd1 _5352_/A sky130_fd_sc_hd__a21o_1
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5276_ _5276_/A _5386_/A vssd1 vssd1 vccd1 vccd1 _5276_/X sky130_fd_sc_hd__or2_1
X_7015_ _5987_/A _7005_/X _7014_/X _7007_/X vssd1 vssd1 vccd1 vccd1 _7184_/D sky130_fd_sc_hd__o211a_1
X_4227_ _7178_/Q vssd1 vssd1 vccd1 vccd1 hold90/A sky130_fd_sc_hd__buf_2
XFILLER_46_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4158_ _4158_/A _4158_/B vssd1 vssd1 vccd1 vccd1 _4159_/B sky130_fd_sc_hd__nor2_1
XFILLER_55_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7282__75 vssd1 vssd1 vccd1 vccd1 _7282__75/HI _7381_/A sky130_fd_sc_hd__conb_1
X_4089_ _4329_/A vssd1 vssd1 vccd1 vccd1 _5019_/A sky130_fd_sc_hd__buf_2
XFILLER_43_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput13 io_in[21] vssd1 vssd1 vccd1 vccd1 _6886_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_97_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5130_ _5286_/A _5286_/B vssd1 vssd1 vccd1 vccd1 _5135_/A sky130_fd_sc_hd__nor2_1
XFILLER_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5061_ hold84/X vssd1 vssd1 vccd1 vccd1 _7072_/A sky130_fd_sc_hd__inv_2
XFILLER_96_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4012_ _4012_/A _4012_/B _4964_/A vssd1 vssd1 vccd1 vccd1 _4016_/B sky130_fd_sc_hd__or3b_2
XFILLER_65_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5963_ _5963_/A _5963_/B vssd1 vssd1 vccd1 vccd1 _5969_/B sky130_fd_sc_hd__xor2_1
XFILLER_52_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4914_ _5734_/A _4914_/B vssd1 vssd1 vccd1 vccd1 _5630_/A sky130_fd_sc_hd__and2_4
X_5894_ _5894_/A _5894_/B vssd1 vssd1 vccd1 vccd1 _5930_/A sky130_fd_sc_hd__xnor2_1
X_4845_ _5829_/B _6409_/B vssd1 vssd1 vccd1 vccd1 _4847_/B sky130_fd_sc_hd__or2_1
XFILLER_60_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4776_ _4776_/A _4775_/A vssd1 vssd1 vccd1 vccd1 _4776_/X sky130_fd_sc_hd__or2b_1
X_6515_ _6520_/A _6520_/B _6513_/X _6522_/A vssd1 vssd1 vccd1 vccd1 _6515_/X sky130_fd_sc_hd__o211a_1
X_3727_ _3727_/A vssd1 vssd1 vccd1 vccd1 _3727_/Y sky130_fd_sc_hd__inv_2
X_6446_ _6466_/B _6821_/A vssd1 vssd1 vccd1 vccd1 _6448_/A sky130_fd_sc_hd__xnor2_1
X_3658_ _3660_/A vssd1 vssd1 vccd1 vccd1 _3658_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6377_ _6377_/A vssd1 vssd1 vccd1 vccd1 _6378_/B sky130_fd_sc_hd__inv_2
XFILLER_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5328_ _7174_/Q vssd1 vssd1 vccd1 vccd1 _5784_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5259_ _5257_/X _5375_/B hold63/X vssd1 vssd1 vccd1 vccd1 _5259_/X sky130_fd_sc_hd__a21o_1
XFILLER_56_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4630_ _4636_/A _4636_/B _4629_/Y vssd1 vssd1 vccd1 vccd1 _5108_/B sky130_fd_sc_hd__a21o_1
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4561_ _4559_/A _4559_/B _4603_/A vssd1 vssd1 vccd1 vccd1 _4597_/A sky130_fd_sc_hd__a21o_1
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6300_ _6300_/A _6349_/B vssd1 vssd1 vccd1 vccd1 _6305_/A sky130_fd_sc_hd__xor2_2
X_4492_ _4440_/B _4492_/B vssd1 vssd1 vccd1 vccd1 _4493_/B sky130_fd_sc_hd__and2b_1
X_6231_ _6302_/A _6302_/B vssd1 vssd1 vccd1 vccd1 _6233_/A sky130_fd_sc_hd__or2_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ _6528_/A _6162_/B _6162_/C _5801_/A vssd1 vssd1 vccd1 vccd1 _6163_/B sky130_fd_sc_hd__or4b_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5113_ _6845_/A vssd1 vssd1 vccd1 vccd1 _5113_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_97_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ _5862_/A _5862_/B _6092_/Y vssd1 vssd1 vccd1 vccd1 _6189_/B sky130_fd_sc_hd__a21oi_2
XFILLER_84_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5044_ _4388_/A _5042_/X _5043_/X vssd1 vssd1 vccd1 vccd1 _5095_/A sky130_fd_sc_hd__o21a_1
X_7252__45 vssd1 vssd1 vccd1 vccd1 _7252__45/HI _7351_/A sky130_fd_sc_hd__conb_1
XFILLER_25_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6995_ _7007_/A vssd1 vssd1 vccd1 vccd1 _6995_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5946_ _5985_/B _5739_/D _5897_/Y vssd1 vssd1 vccd1 vccd1 _5975_/A sky130_fd_sc_hd__o21ai_2
XFILLER_80_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5877_ _5630_/A _4916_/B _5911_/B _5876_/B _5876_/A vssd1 vssd1 vccd1 vccd1 _5879_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_21_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4828_ _4869_/A _4869_/B _4827_/Y vssd1 vssd1 vccd1 vccd1 _4830_/B sky130_fd_sc_hd__o21a_1
X_4759_ _4759_/A _4759_/B vssd1 vssd1 vccd1 vccd1 _4814_/A sky130_fd_sc_hd__xor2_1
X_6429_ _6466_/A vssd1 vssd1 vccd1 vccd1 _6588_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_88_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_66_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3992_ _4014_/B vssd1 vssd1 vccd1 vccd1 _3992_/Y sky130_fd_sc_hd__inv_2
X_6780_ _6792_/A _6792_/B vssd1 vssd1 vccd1 vccd1 _6793_/B sky130_fd_sc_hd__xor2_1
X_5800_ _6085_/B _5800_/B vssd1 vssd1 vccd1 vccd1 _5810_/A sky130_fd_sc_hd__xnor2_2
X_5731_ _5730_/B _5731_/B vssd1 vssd1 vccd1 vccd1 _5731_/X sky130_fd_sc_hd__and2b_1
XFILLER_50_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5662_ _6014_/A _6014_/B _6020_/A vssd1 vssd1 vccd1 vccd1 _5663_/B sky130_fd_sc_hd__o21a_1
X_4613_ _4613_/A _4694_/B _4613_/C vssd1 vssd1 vccd1 vccd1 _4614_/S sky130_fd_sc_hd__or3_1
X_7401_ _7401_/A _3695_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[5] sky130_fd_sc_hd__ebufn_8
X_5593_ hold63/X hold13/X _5590_/X _5592_/Y _6907_/A vssd1 vssd1 vccd1 vccd1 hold76/A
+ sky130_fd_sc_hd__a221oi_1
XFILLER_30_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4544_ _4641_/A _4642_/A _4641_/B _4542_/A vssd1 vssd1 vccd1 vccd1 _4545_/A sky130_fd_sc_hd__o31a_1
X_7332_ _7332_/A _3612_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[6] sky130_fd_sc_hd__ebufn_8
X_4475_ _4488_/A _4488_/B vssd1 vssd1 vccd1 vccd1 _4562_/A sky130_fd_sc_hd__xor2_1
X_6214_ _4375_/B _4298_/Y _6039_/B vssd1 vssd1 vccd1 vccd1 _6215_/B sky130_fd_sc_hd__o21a_1
X_7194_ _7221_/CLK _7194_/D vssd1 vssd1 vccd1 vccd1 _7194_/Q sky130_fd_sc_hd__dfxtp_2
X_6145_ _6145_/A _6145_/B vssd1 vssd1 vccd1 vccd1 _6146_/B sky130_fd_sc_hd__xor2_4
XFILLER_38_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6076_ _6076_/A _6076_/B _6076_/C vssd1 vssd1 vccd1 vccd1 _6078_/A sky130_fd_sc_hd__nor3_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5027_ _6956_/A _6470_/A _5024_/X vssd1 vssd1 vccd1 vccd1 _5028_/B sky130_fd_sc_hd__a21o_1
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6978_ _6978_/A _6983_/B vssd1 vssd1 vccd1 vccd1 _6978_/Y sky130_fd_sc_hd__nand2_1
X_5929_ _5941_/A _5941_/B _5928_/X vssd1 vssd1 vccd1 vccd1 _5930_/B sky130_fd_sc_hd__a21oi_1
XFILLER_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4260_ _4260_/A _4260_/B _4260_/C vssd1 vssd1 vccd1 vccd1 _4260_/X sky130_fd_sc_hd__or3_1
X_4191_ _7210_/Q _7209_/Q vssd1 vssd1 vccd1 vccd1 _4540_/B sky130_fd_sc_hd__and2_1
XFILLER_79_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6901_ hold19/X _6892_/X _6894_/X hold17/X vssd1 vssd1 vccd1 vccd1 _6901_/X sky130_fd_sc_hd__a22o_1
XFILLER_35_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6832_ _6850_/A _6850_/B vssd1 vssd1 vccd1 vccd1 _6835_/A sky130_fd_sc_hd__xor2_1
XFILLER_35_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3975_ _5029_/A _3975_/B vssd1 vssd1 vccd1 vccd1 _3980_/A sky130_fd_sc_hd__nor2_2
XFILLER_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6763_ _6763_/A _6763_/B vssd1 vssd1 vccd1 vccd1 _6763_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6694_ _6971_/A _6926_/A vssd1 vssd1 vccd1 vccd1 _6694_/X sky130_fd_sc_hd__and2b_1
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5714_ _5714_/A _5714_/B vssd1 vssd1 vccd1 vccd1 _5759_/A sky130_fd_sc_hd__xor2_2
X_5645_ _6674_/A vssd1 vssd1 vccd1 vccd1 _5936_/A sky130_fd_sc_hd__inv_2
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5576_ _5574_/X _5575_/Y _5567_/B _5570_/A vssd1 vssd1 vccd1 vccd1 _5590_/A sky130_fd_sc_hd__a31o_1
X_4527_ _4527_/A _4527_/B vssd1 vssd1 vccd1 vccd1 _4529_/B sky130_fd_sc_hd__xnor2_1
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4458_ _6120_/B _4458_/B vssd1 vssd1 vccd1 vccd1 _4470_/B sky130_fd_sc_hd__xnor2_1
XFILLER_77_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7177_ _7225_/CLK _7177_/D vssd1 vssd1 vccd1 vccd1 _7177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4389_ _4389_/A _4389_/B vssd1 vssd1 vccd1 vccd1 _4390_/B sky130_fd_sc_hd__xnor2_2
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6128_ _6116_/B _6128_/B vssd1 vssd1 vccd1 vccd1 _6128_/X sky130_fd_sc_hd__and2b_1
XFILLER_85_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6059_ _6171_/A _6171_/B vssd1 vssd1 vccd1 vccd1 _6079_/A sky130_fd_sc_hd__xnor2_2
XFILLER_45_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7288__81 vssd1 vssd1 vccd1 vccd1 _7288__81/HI _7396_/A sky130_fd_sc_hd__conb_1
XFILLER_1_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3760_ _5198_/B _5625_/B vssd1 vssd1 vccd1 vccd1 _3761_/C sky130_fd_sc_hd__nand2_1
XFILLER_32_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3691_ _3691_/A vssd1 vssd1 vccd1 vccd1 _3691_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5430_ _5430_/A vssd1 vssd1 vccd1 vccd1 _6575_/A sky130_fd_sc_hd__clkbuf_4
X_5361_ _5361_/A _5361_/B vssd1 vssd1 vccd1 vccd1 _5361_/Y sky130_fd_sc_hd__nand2_1
X_4312_ _4460_/A _5871_/A vssd1 vssd1 vccd1 vccd1 _4452_/B sky130_fd_sc_hd__xnor2_1
X_7100_ _7078_/A _7088_/X hold81/X _7099_/X vssd1 vssd1 vccd1 vccd1 _7216_/D sky130_fd_sc_hd__o211a_1
X_5292_ _5292_/A _6945_/A vssd1 vssd1 vccd1 vccd1 _5293_/B sky130_fd_sc_hd__nand2_1
X_4243_ _4243_/A _4243_/B vssd1 vssd1 vccd1 vccd1 _4497_/A sky130_fd_sc_hd__xnor2_4
XFILLER_87_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7031_ _7009_/A _7018_/X _7030_/X _7021_/X vssd1 vssd1 vccd1 vccd1 _7190_/D sky130_fd_sc_hd__o211a_1
X_4174_ _4173_/B _4174_/B vssd1 vssd1 vccd1 vccd1 _4174_/X sky130_fd_sc_hd__and2b_1
XFILLER_67_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6815_ _6815_/A vssd1 vssd1 vccd1 vccd1 _6816_/B sky130_fd_sc_hd__inv_2
XFILLER_11_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6746_ _6585_/A _6585_/B _6745_/X vssd1 vssd1 vccd1 vccd1 _6747_/B sky130_fd_sc_hd__o21a_1
X_3958_ _6110_/A vssd1 vssd1 vccd1 vccd1 _6941_/A sky130_fd_sc_hd__inv_2
X_6677_ _6677_/A _6677_/B vssd1 vssd1 vccd1 vccd1 _6682_/A sky130_fd_sc_hd__nand2_1
X_3889_ _3889_/A _3889_/B _3889_/C vssd1 vssd1 vccd1 vccd1 _3890_/B sky130_fd_sc_hd__or3_1
X_5628_ _6659_/A _5983_/A vssd1 vssd1 vccd1 vccd1 _5628_/Y sky130_fd_sc_hd__nor2_1
X_5559_ _5559_/A _5578_/B vssd1 vssd1 vccd1 vccd1 _5563_/A sky130_fd_sc_hd__xor2_1
XFILLER_58_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_1_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7183_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_42_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4930_ _4924_/X _4926_/Y _4929_/Y _4931_/B _4931_/A vssd1 vssd1 vccd1 vccd1 _4934_/A
+ sky130_fd_sc_hd__a32o_1
X_4861_ _4878_/A _4861_/B vssd1 vssd1 vccd1 vccd1 _4862_/B sky130_fd_sc_hd__and2_1
XFILLER_17_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3812_ _7186_/Q vssd1 vssd1 vccd1 vccd1 _5667_/B sky130_fd_sc_hd__buf_2
X_6600_ _6971_/A _6600_/B vssd1 vssd1 vccd1 vccd1 _6601_/B sky130_fd_sc_hd__nand2_1
X_4792_ _4864_/A _4864_/B vssd1 vssd1 vccd1 vccd1 _4865_/A sky130_fd_sc_hd__nand2_1
XANTENNA_27 _7063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_38 _7117_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_16 _6073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_49 _7106_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3743_ _6907_/A vssd1 vssd1 vccd1 vccd1 _7020_/A sky130_fd_sc_hd__clkinv_2
X_6531_ _6531_/A _6531_/B vssd1 vssd1 vccd1 vccd1 _6533_/B sky130_fd_sc_hd__xnor2_1
X_6462_ _6730_/A _6462_/B vssd1 vssd1 vccd1 vccd1 _6724_/A sky130_fd_sc_hd__nand2_2
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3674_ _3678_/A vssd1 vssd1 vccd1 vccd1 _3674_/Y sky130_fd_sc_hd__inv_2
X_6393_ _6387_/B _6393_/B vssd1 vssd1 vccd1 vccd1 _6393_/X sky130_fd_sc_hd__and2b_1
X_5413_ _5413_/A _5413_/B vssd1 vssd1 vccd1 vccd1 _5414_/B sky130_fd_sc_hd__or2_1
X_5344_ _6270_/A vssd1 vssd1 vccd1 vccd1 _5450_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5275_ _5275_/A _7055_/A vssd1 vssd1 vccd1 vccd1 _5386_/A sky130_fd_sc_hd__nand2_1
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7014_ _7014_/A _7025_/B vssd1 vssd1 vccd1 vccd1 _7014_/X sky130_fd_sc_hd__or2_1
X_4226_ _6722_/A _4226_/B vssd1 vssd1 vccd1 vccd1 _4293_/A sky130_fd_sc_hd__xnor2_2
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4157_ _4157_/A _4157_/B _4157_/C vssd1 vssd1 vccd1 vccd1 _4158_/B sky130_fd_sc_hd__and3_1
X_4088_ _7163_/Q vssd1 vssd1 vccd1 vccd1 _4329_/A sky130_fd_sc_hd__buf_2
XFILLER_83_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6729_ _6767_/A _6729_/B vssd1 vssd1 vccd1 vccd1 _6730_/C sky130_fd_sc_hd__nand2_1
XFILLER_11_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7258__51 vssd1 vssd1 vccd1 vccd1 _7258__51/HI _7357_/A sky130_fd_sc_hd__conb_1
XFILLER_100_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput14 io_in[22] vssd1 vssd1 vccd1 vccd1 _6886_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5060_ hold85/X vssd1 vssd1 vccd1 vccd1 hold84/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4011_ _4011_/A _4011_/B vssd1 vssd1 vccd1 vccd1 _4964_/A sky130_fd_sc_hd__nor2_2
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5962_ _6007_/A _5962_/B vssd1 vssd1 vccd1 vccd1 _5969_/A sky130_fd_sc_hd__nand2_1
XFILLER_65_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4913_ _5987_/A _4910_/X _4912_/X vssd1 vssd1 vccd1 vccd1 _4913_/X sky130_fd_sc_hd__o21a_1
XFILLER_52_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5893_ _5893_/A _5893_/B vssd1 vssd1 vccd1 vccd1 _5934_/A sky130_fd_sc_hd__xnor2_1
X_4844_ _4844_/A vssd1 vssd1 vccd1 vccd1 _6409_/B sky130_fd_sc_hd__buf_2
XFILLER_21_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4775_ _4775_/A _4776_/A vssd1 vssd1 vccd1 vccd1 _4814_/B sky130_fd_sc_hd__xnor2_1
X_6514_ _6514_/A _6514_/B vssd1 vssd1 vccd1 vccd1 _6522_/A sky130_fd_sc_hd__xor2_2
X_3726_ _3727_/A vssd1 vssd1 vccd1 vccd1 _3726_/Y sky130_fd_sc_hd__inv_2
X_6445_ _7159_/Q _6445_/B vssd1 vssd1 vccd1 vccd1 _6821_/A sky130_fd_sc_hd__xnor2_4
X_3657_ _3660_/A vssd1 vssd1 vccd1 vccd1 _3657_/Y sky130_fd_sc_hd__inv_2
X_6376_ _6874_/A _6375_/B _6375_/Y vssd1 vssd1 vccd1 vccd1 _6377_/A sky130_fd_sc_hd__o21a_1
XFILLER_88_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5327_ _5446_/A _5446_/B vssd1 vssd1 vccd1 vccd1 _5340_/A sky130_fd_sc_hd__nand2_1
XFILLER_75_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5258_ _5257_/A _5257_/B _5257_/C vssd1 vssd1 vccd1 vccd1 _5375_/B sky130_fd_sc_hd__o21ai_1
X_4209_ hold94/A _6507_/A vssd1 vssd1 vccd1 vccd1 _4210_/B sky130_fd_sc_hd__nor2_1
XFILLER_68_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5189_ _3783_/A _5048_/A _5190_/B _5054_/B _5054_/A vssd1 vssd1 vccd1 vccd1 _5202_/A
+ sky130_fd_sc_hd__a32o_2
XFILLER_73_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4560_ _4602_/B _4560_/B vssd1 vssd1 vccd1 vccd1 _4603_/A sky130_fd_sc_hd__and2b_1
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4491_ _4491_/A _4491_/B vssd1 vssd1 vccd1 vccd1 _4520_/A sky130_fd_sc_hd__xnor2_4
X_6230_ _6230_/A _6230_/B vssd1 vssd1 vccd1 vccd1 _6302_/B sky130_fd_sc_hd__or2_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6161_ _5801_/A _6158_/Y _6162_/B vssd1 vssd1 vccd1 vccd1 _6234_/A sky130_fd_sc_hd__a21bo_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ _5111_/A _5111_/B _5111_/C vssd1 vssd1 vccd1 vccd1 _5257_/B sky130_fd_sc_hd__a21oi_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6092_ _6092_/A _6092_/B vssd1 vssd1 vccd1 vccd1 _6092_/Y sky130_fd_sc_hd__nor2_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5043_ _5043_/A _5043_/B vssd1 vssd1 vccd1 vccd1 _5043_/X sky130_fd_sc_hd__or2_1
XFILLER_38_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6994_ _6994_/A _7006_/B vssd1 vssd1 vccd1 vccd1 _6994_/Y sky130_fd_sc_hd__nand2_1
X_5945_ _5945_/A _5945_/B vssd1 vssd1 vccd1 vccd1 _5978_/A sky130_fd_sc_hd__or2_1
X_5876_ _5876_/A _5876_/B vssd1 vssd1 vccd1 vccd1 _5911_/B sky130_fd_sc_hd__xnor2_2
XFILLER_40_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4827_ _4827_/A _4827_/B vssd1 vssd1 vccd1 vccd1 _4827_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4758_ _4758_/A _4758_/B vssd1 vssd1 vccd1 vccd1 _4778_/A sky130_fd_sc_hd__xnor2_1
X_3709_ _3709_/A vssd1 vssd1 vccd1 vccd1 _3709_/Y sky130_fd_sc_hd__inv_2
X_4689_ _4689_/A _4689_/B vssd1 vssd1 vccd1 vccd1 _4756_/A sky130_fd_sc_hd__xor2_1
X_6428_ _6720_/A _6428_/B vssd1 vssd1 vccd1 vccd1 _6536_/A sky130_fd_sc_hd__or2_1
X_6359_ _6359_/A _6359_/B vssd1 vssd1 vccd1 vccd1 _6359_/X sky130_fd_sc_hd__xor2_1
XFILLER_88_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7228__21 vssd1 vssd1 vccd1 vccd1 _7228__21/HI _7327_/A sky130_fd_sc_hd__conb_1
XFILLER_48_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_74_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3991_ _4694_/A _4172_/B _3990_/X vssd1 vssd1 vccd1 vccd1 _4014_/B sky130_fd_sc_hd__a21oi_2
XFILLER_74_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5730_ _5731_/B _5730_/B vssd1 vssd1 vccd1 vccd1 _5759_/B sky130_fd_sc_hd__xnor2_2
X_5661_ _6022_/A _6483_/B vssd1 vssd1 vccd1 vccd1 _6020_/B sky130_fd_sc_hd__xor2_4
X_7400_ _7400_/A _3694_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[4] sky130_fd_sc_hd__ebufn_8
X_4612_ _5722_/A vssd1 vssd1 vccd1 vccd1 _7023_/A sky130_fd_sc_hd__buf_2
X_5592_ _5590_/A _5590_/B _6879_/A vssd1 vssd1 vccd1 vccd1 _5592_/Y sky130_fd_sc_hd__a21oi_1
X_4543_ _4543_/A _4543_/B vssd1 vssd1 vccd1 vccd1 _4641_/B sky130_fd_sc_hd__nor2_1
X_7331_ _7331_/A _3742_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[5] sky130_fd_sc_hd__ebufn_8
X_4474_ _4474_/A _4586_/A vssd1 vssd1 vccd1 vccd1 _4488_/B sky130_fd_sc_hd__nor2_1
X_6213_ _6213_/A _6213_/B vssd1 vssd1 vccd1 vccd1 _6215_/A sky130_fd_sc_hd__xnor2_2
X_7193_ _7221_/CLK _7193_/D vssd1 vssd1 vccd1 vccd1 _7193_/Q sky130_fd_sc_hd__dfxtp_1
X_6144_ _7003_/A _6329_/A _6143_/X vssd1 vssd1 vccd1 vccd1 _6145_/B sky130_fd_sc_hd__a21oi_2
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6075_ _6075_/A _6075_/B vssd1 vssd1 vccd1 vccd1 _6076_/C sky130_fd_sc_hd__xnor2_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5026_ _5026_/A vssd1 vssd1 vccd1 vccd1 _6956_/A sky130_fd_sc_hd__clkbuf_4
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6977_ _6977_/A vssd1 vssd1 vccd1 vccd1 _6977_/X sky130_fd_sc_hd__clkbuf_2
X_5928_ _5927_/B _5928_/B vssd1 vssd1 vccd1 vccd1 _5928_/X sky130_fd_sc_hd__and2b_1
X_5859_ _5859_/A _5859_/B _5859_/C vssd1 vssd1 vccd1 vccd1 _5860_/B sky130_fd_sc_hd__nor3_1
XFILLER_5_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4190_ _7210_/Q _7209_/Q vssd1 vssd1 vccd1 vccd1 _4726_/B sky130_fd_sc_hd__or2_1
XFILLER_94_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6900_ _6906_/A hold34/X vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__nor2_1
XFILLER_35_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6831_ _6831_/A _6849_/B vssd1 vssd1 vccd1 vccd1 _6850_/B sky130_fd_sc_hd__xor2_1
XFILLER_35_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3974_ hold96/A _3974_/B vssd1 vssd1 vccd1 vccd1 _3975_/B sky130_fd_sc_hd__and2_1
X_6762_ _4308_/B _6761_/B _6761_/Y vssd1 vssd1 vccd1 vccd1 _6773_/A sky130_fd_sc_hd__a21o_1
XFILLER_50_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6693_ _6693_/A _6693_/B vssd1 vssd1 vccd1 vccd1 _6693_/Y sky130_fd_sc_hd__nand2_1
X_5713_ _5762_/A _4321_/A _5718_/A vssd1 vssd1 vccd1 vccd1 _5714_/B sky130_fd_sc_hd__mux2_1
X_5644_ _5644_/A vssd1 vssd1 vccd1 vccd1 _6674_/A sky130_fd_sc_hd__clkbuf_2
X_5575_ _5575_/A _5575_/B vssd1 vssd1 vccd1 vccd1 _5575_/Y sky130_fd_sc_hd__nand2_1
X_4526_ _4533_/A _4526_/B _4873_/A vssd1 vssd1 vccd1 vccd1 _4611_/A sky130_fd_sc_hd__and3_1
X_4457_ _4472_/A _4472_/B vssd1 vssd1 vccd1 vccd1 _4474_/A sky130_fd_sc_hd__and2b_1
X_7176_ _7225_/CLK _7176_/D vssd1 vssd1 vccd1 vccd1 _7176_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6127_ _6270_/A _6127_/B vssd1 vssd1 vccd1 vccd1 _6198_/A sky130_fd_sc_hd__xnor2_2
X_4388_ _4388_/A _4388_/B vssd1 vssd1 vccd1 vccd1 _4389_/B sky130_fd_sc_hd__xnor2_4
XFILLER_100_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6058_ _6056_/Y _5748_/B _6057_/Y vssd1 vssd1 vccd1 vccd1 _6171_/B sky130_fd_sc_hd__a21oi_2
XFILLER_45_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5009_ _5690_/A _5784_/B vssd1 vssd1 vccd1 vccd1 _5228_/B sky130_fd_sc_hd__xor2_2
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3690_ _3691_/A vssd1 vssd1 vccd1 vccd1 _3690_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5360_ _5360_/A _5360_/B vssd1 vssd1 vccd1 vccd1 _5464_/A sky130_fd_sc_hd__xnor2_1
XFILLER_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4311_ _4311_/A vssd1 vssd1 vccd1 vccd1 _5871_/A sky130_fd_sc_hd__clkbuf_2
X_5291_ _6464_/A vssd1 vssd1 vccd1 vccd1 _6945_/A sky130_fd_sc_hd__clkbuf_4
X_4242_ _4260_/A _4260_/B vssd1 vssd1 vccd1 vccd1 _4259_/A sky130_fd_sc_hd__nor2_1
X_7030_ _7053_/A _7038_/B vssd1 vssd1 vccd1 vccd1 _7030_/X sky130_fd_sc_hd__or2_1
X_4173_ _4174_/B _4173_/B vssd1 vssd1 vccd1 vccd1 _4247_/A sky130_fd_sc_hd__xnor2_2
XFILLER_95_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6814_ _6814_/A _6814_/B _6814_/C vssd1 vssd1 vccd1 vccd1 _6815_/A sky130_fd_sc_hd__nand3_1
X_3957_ _6484_/A vssd1 vssd1 vccd1 vccd1 _6110_/A sky130_fd_sc_hd__clkbuf_2
X_6745_ _6745_/A _6583_/A vssd1 vssd1 vccd1 vccd1 _6745_/X sky130_fd_sc_hd__or2b_1
XFILLER_50_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6676_ _6676_/A vssd1 vssd1 vccd1 vccd1 _6677_/B sky130_fd_sc_hd__inv_2
X_3888_ _3889_/A _3889_/B _3889_/C vssd1 vssd1 vccd1 vccd1 _4992_/A sky130_fd_sc_hd__o21ai_1
X_5627_ _5736_/C _5627_/B vssd1 vssd1 vccd1 vccd1 _5983_/A sky130_fd_sc_hd__nand2_2
X_5558_ _5558_/A _5558_/B vssd1 vssd1 vccd1 vccd1 _5578_/B sky130_fd_sc_hd__nand2_1
X_4509_ _4638_/B _4613_/C _4507_/A _4503_/Y _4508_/Y vssd1 vssd1 vccd1 vccd1 _4511_/B
+ sky130_fd_sc_hd__o41a_1
X_5489_ _5490_/A _5490_/B _5490_/C vssd1 vssd1 vccd1 vccd1 _5551_/A sky130_fd_sc_hd__o21ai_1
X_7159_ _7172_/CLK _7159_/D vssd1 vssd1 vccd1 vccd1 _7159_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4860_ _4878_/A _4861_/B vssd1 vssd1 vccd1 vccd1 _4867_/A sky130_fd_sc_hd__nor2_1
X_3811_ _3811_/A _4339_/B vssd1 vssd1 vccd1 vccd1 _4632_/A sky130_fd_sc_hd__nor2_2
XFILLER_60_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_28 _7045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4791_ _4791_/A _4791_/B vssd1 vssd1 vccd1 vccd1 _4864_/B sky130_fd_sc_hd__nor2_1
XANTENNA_17 _6111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_39 _7117_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6530_ _6539_/A _6539_/B vssd1 vssd1 vccd1 vccd1 _6540_/A sky130_fd_sc_hd__nor2_1
XFILLER_32_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3742_ _3742_/A vssd1 vssd1 vccd1 vccd1 _3742_/Y sky130_fd_sc_hd__inv_2
X_6461_ _6461_/A _6460_/A vssd1 vssd1 vccd1 vccd1 _6462_/B sky130_fd_sc_hd__or2b_1
X_3673_ _3679_/A vssd1 vssd1 vccd1 vccd1 _3678_/A sky130_fd_sc_hd__buf_2
XFILLER_9_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6392_ _6261_/X _6390_/X _6391_/X _6196_/X vssd1 vssd1 vccd1 vccd1 _7134_/D sky130_fd_sc_hd__o211a_1
X_5412_ _6270_/A _5412_/B _5412_/C vssd1 vssd1 vccd1 vccd1 _5413_/B sky130_fd_sc_hd__and3_1
X_5343_ _5381_/A _5381_/B vssd1 vssd1 vccd1 vccd1 _5420_/A sky130_fd_sc_hd__xnor2_1
X_5274_ _5274_/A vssd1 vssd1 vccd1 vccd1 _5391_/B sky130_fd_sc_hd__buf_2
X_7013_ _7063_/A vssd1 vssd1 vccd1 vccd1 _7025_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4225_ _4225_/A _4225_/B vssd1 vssd1 vccd1 vccd1 _4226_/B sky130_fd_sc_hd__xnor2_2
X_4156_ _4157_/A _4157_/B _4157_/C vssd1 vssd1 vccd1 vccd1 _4158_/A sky130_fd_sc_hd__a21oi_1
XFILLER_28_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4087_ _4572_/A vssd1 vssd1 vccd1 vccd1 _4573_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4989_ _4989_/A _4989_/B vssd1 vssd1 vccd1 vccd1 _4990_/B sky130_fd_sc_hd__nor2_1
X_6728_ _6728_/A _6727_/B vssd1 vssd1 vccd1 vccd1 _6729_/B sky130_fd_sc_hd__or2b_1
X_6659_ _6659_/A vssd1 vssd1 vccd1 vccd1 _6659_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7273__66 vssd1 vssd1 vccd1 vccd1 _7273__66/HI _7372_/A sky130_fd_sc_hd__conb_1
XFILLER_46_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput15 io_in[23] vssd1 vssd1 vccd1 vccd1 _6886_/D sky130_fd_sc_hd__buf_2
XFILLER_10_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7323__116 vssd1 vssd1 vccd1 vccd1 _7323__116/HI _7431_/A sky130_fd_sc_hd__conb_1
X_4010_ _3844_/X _4009_/B _4506_/C vssd1 vssd1 vccd1 vccd1 _4012_/B sky130_fd_sc_hd__a21oi_1
X_5961_ _6693_/A _4328_/B _5954_/A vssd1 vssd1 vccd1 vccd1 _5962_/B sky130_fd_sc_hd__a21o_1
X_4912_ _5880_/B _4910_/X _4911_/X _4899_/B vssd1 vssd1 vccd1 vccd1 _4912_/X sky130_fd_sc_hd__a22o_1
X_5892_ _6097_/A _6097_/B vssd1 vssd1 vccd1 vccd1 _5893_/B sky130_fd_sc_hd__xor2_2
X_4843_ _6502_/B vssd1 vssd1 vccd1 vccd1 _5829_/B sky130_fd_sc_hd__buf_2
X_4774_ _4772_/A _4772_/B _4817_/A vssd1 vssd1 vccd1 vccd1 _4776_/A sky130_fd_sc_hd__a21oi_2
X_6513_ _6520_/A _6520_/B _6512_/X vssd1 vssd1 vccd1 vccd1 _6513_/X sky130_fd_sc_hd__a21o_1
X_3725_ _3727_/A vssd1 vssd1 vccd1 vccd1 _3725_/Y sky130_fd_sc_hd__inv_2
X_6444_ _6481_/A _6481_/B _6443_/Y vssd1 vssd1 vccd1 vccd1 _6460_/A sky130_fd_sc_hd__a21oi_1
X_3656_ _3660_/A vssd1 vssd1 vccd1 vccd1 _3656_/Y sky130_fd_sc_hd__inv_2
X_6375_ _6986_/A _6375_/B vssd1 vssd1 vccd1 vccd1 _6375_/Y sky130_fd_sc_hd__nand2_1
XFILLER_88_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5326_ _5181_/A _5181_/B _5325_/X vssd1 vssd1 vccd1 vccd1 _5358_/A sky130_fd_sc_hd__a21o_1
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5257_ _5257_/A _5257_/B _5257_/C vssd1 vssd1 vccd1 vccd1 _5257_/X sky130_fd_sc_hd__or3_1
X_4208_ _4208_/A _4429_/A _6479_/B vssd1 vssd1 vccd1 vccd1 _4422_/A sky130_fd_sc_hd__and3_1
XFILLER_68_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5188_ _5341_/A _5341_/B vssd1 vssd1 vccd1 vccd1 _5219_/A sky130_fd_sc_hd__nand2_1
X_4139_ _5168_/A _6617_/A vssd1 vssd1 vccd1 vccd1 _4139_/Y sky130_fd_sc_hd__nand2_1
XFILLER_71_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4490_ _4523_/A _4523_/B vssd1 vssd1 vccd1 vccd1 _4599_/A sky130_fd_sc_hd__xor2_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6160_ _6160_/A _6160_/B vssd1 vssd1 vccd1 vccd1 _6162_/B sky130_fd_sc_hd__xnor2_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5111_ _5111_/A _5111_/B _5111_/C vssd1 vssd1 vccd1 vccd1 _5111_/X sky130_fd_sc_hd__and3_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _6091_/A _6091_/B vssd1 vssd1 vccd1 vccd1 _6189_/A sky130_fd_sc_hd__xnor2_4
XFILLER_84_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _5043_/A _5043_/B vssd1 vssd1 vccd1 vccd1 _5042_/X sky130_fd_sc_hd__and2_1
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6993_ _7045_/A vssd1 vssd1 vccd1 vccd1 _6993_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_25_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5944_ _6994_/A _5944_/B vssd1 vssd1 vccd1 vccd1 _5945_/B sky130_fd_sc_hd__and2_1
X_5875_ hold89/A _5912_/B _5912_/A vssd1 vssd1 vccd1 vccd1 _5876_/B sky130_fd_sc_hd__a21boi_2
XFILLER_21_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4826_ _4827_/A _4827_/B vssd1 vssd1 vccd1 vccd1 _4869_/B sky130_fd_sc_hd__xnor2_2
XFILLER_21_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4757_ _4757_/A _4757_/B vssd1 vssd1 vccd1 vccd1 _4812_/A sky130_fd_sc_hd__xor2_1
X_4688_ _4688_/A _4688_/B vssd1 vssd1 vccd1 vccd1 _4714_/A sky130_fd_sc_hd__xnor2_1
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3708_ _3709_/A vssd1 vssd1 vccd1 vccd1 _3708_/Y sky130_fd_sc_hd__inv_2
X_3639_ _3641_/A vssd1 vssd1 vccd1 vccd1 _3639_/Y sky130_fd_sc_hd__inv_2
X_6427_ _6975_/A _6552_/A vssd1 vssd1 vccd1 vccd1 _6428_/B sky130_fd_sc_hd__and2_1
X_6358_ _6319_/A _6319_/B _6357_/X vssd1 vssd1 vccd1 vccd1 _6359_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5309_ _6034_/A vssd1 vssd1 vccd1 vccd1 _6270_/A sky130_fd_sc_hd__buf_2
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6289_ _6966_/A _6289_/B vssd1 vssd1 vccd1 vccd1 _6290_/C sky130_fd_sc_hd__xnor2_1
XFILLER_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7243__36 vssd1 vssd1 vccd1 vccd1 _7243__36/HI _7342_/A sky130_fd_sc_hd__conb_1
XFILLER_16_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_94_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3990_ _4412_/B _4527_/A vssd1 vssd1 vccd1 vccd1 _3990_/X sky130_fd_sc_hd__and2_1
XFILLER_62_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5660_ _5682_/A _5682_/B vssd1 vssd1 vccd1 vccd1 _5683_/A sky130_fd_sc_hd__nand2_2
XFILLER_30_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4611_ _4611_/A _4611_/B vssd1 vssd1 vccd1 vccd1 _4693_/A sky130_fd_sc_hd__or2_2
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5591_ hold74/X vssd1 vssd1 vccd1 vccd1 _6879_/A sky130_fd_sc_hd__buf_2
XFILLER_30_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4542_ _4542_/A _4542_/B vssd1 vssd1 vccd1 vccd1 _4642_/A sky130_fd_sc_hd__nand2_1
X_7330_ _7330_/A _3741_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[4] sky130_fd_sc_hd__ebufn_8
X_4473_ _4564_/A _4564_/B _4564_/C vssd1 vssd1 vccd1 vccd1 _4586_/A sky130_fd_sc_hd__o21a_1
XFILLER_89_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6212_ _6212_/A _6262_/B vssd1 vssd1 vccd1 vccd1 _6213_/B sky130_fd_sc_hd__xor2_2
X_7192_ _7221_/CLK _7192_/D vssd1 vssd1 vccd1 vccd1 _7192_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_97_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6143_ _6141_/X _6142_/X _6329_/A vssd1 vssd1 vccd1 vccd1 _6143_/X sky130_fd_sc_hd__o21ba_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6074_ _6074_/A _6167_/B vssd1 vssd1 vccd1 vccd1 _6075_/B sky130_fd_sc_hd__nand2_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5025_ _5640_/A _6464_/A _5024_/X vssd1 vssd1 vccd1 vccd1 _5171_/B sky130_fd_sc_hd__or3b_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6976_ _6954_/A _6964_/X _6975_/X _6967_/X vssd1 vssd1 vccd1 vccd1 _7170_/D sky130_fd_sc_hd__o211a_1
XFILLER_26_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5927_ _5928_/B _5927_/B vssd1 vssd1 vccd1 vccd1 _5941_/B sky130_fd_sc_hd__xnor2_1
XFILLER_34_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5858_ _5859_/A _5859_/B _5859_/C vssd1 vssd1 vccd1 vccd1 _5860_/A sky130_fd_sc_hd__o21a_1
X_4809_ _4809_/A _4810_/A vssd1 vssd1 vccd1 vccd1 _4813_/B sky130_fd_sc_hd__xor2_1
X_5789_ _5789_/A _6065_/A vssd1 vssd1 vccd1 vccd1 _5792_/A sky130_fd_sc_hd__xnor2_1
XFILLER_5_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6830_ _6805_/A _6805_/B _6829_/Y vssd1 vssd1 vccd1 vccd1 _6849_/B sky130_fd_sc_hd__o21ai_1
XFILLER_90_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6761_ _6956_/A _6761_/B vssd1 vssd1 vccd1 vccd1 _6761_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5712_ _5717_/A _6137_/B vssd1 vssd1 vccd1 vccd1 _5718_/A sky130_fd_sc_hd__nand2_2
X_3973_ hold96/A _3974_/B vssd1 vssd1 vccd1 vccd1 _5029_/A sky130_fd_sc_hd__nor2_2
XFILLER_50_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6692_ _6950_/A _6693_/B _6690_/B vssd1 vssd1 vccd1 vccd1 _6692_/X sky130_fd_sc_hd__a21bo_1
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5643_ _5643_/A _5643_/B vssd1 vssd1 vccd1 vccd1 _5647_/A sky130_fd_sc_hd__nand2_1
X_5574_ _5575_/A _5575_/B vssd1 vssd1 vccd1 vccd1 _5574_/X sky130_fd_sc_hd__or2_1
X_4525_ _4525_/A _5104_/A vssd1 vssd1 vccd1 vccd1 _5108_/A sky130_fd_sc_hd__xnor2_1
X_4456_ _4456_/A _4456_/B vssd1 vssd1 vccd1 vccd1 _4472_/B sky130_fd_sc_hd__xnor2_1
X_7175_ _7183_/CLK _7175_/D vssd1 vssd1 vccd1 vccd1 _7175_/Q sky130_fd_sc_hd__dfxtp_1
X_4387_ _5043_/A _5043_/B vssd1 vssd1 vccd1 vccd1 _4388_/B sky130_fd_sc_hd__xor2_2
XFILLER_100_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6126_ _6210_/A _6210_/B vssd1 vssd1 vccd1 vccd1 _6127_/B sky130_fd_sc_hd__xor2_2
XFILLER_98_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6057_ _6057_/A _6057_/B vssd1 vssd1 vccd1 vccd1 _6057_/Y sky130_fd_sc_hd__nor2_1
XFILLER_85_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5008_ _7183_/Q vssd1 vssd1 vccd1 vccd1 _5690_/A sky130_fd_sc_hd__buf_2
XFILLER_26_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6959_ _7114_/B vssd1 vssd1 vccd1 vccd1 _6975_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4310_ _4310_/A _4745_/B vssd1 vssd1 vccd1 vccd1 _4311_/A sky130_fd_sc_hd__and2_1
X_5290_ _5290_/A _5290_/B vssd1 vssd1 vccd1 vccd1 _5294_/A sky130_fd_sc_hd__nor2_1
X_7279__72 vssd1 vssd1 vccd1 vccd1 _7279__72/HI _7378_/A sky130_fd_sc_hd__conb_1
XFILLER_99_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4241_ _4240_/A _4240_/C _4240_/B vssd1 vssd1 vccd1 vccd1 _4260_/B sky130_fd_sc_hd__a21oi_1
XFILLER_95_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4172_ _4694_/A _4172_/B vssd1 vssd1 vccd1 vccd1 _4173_/B sky130_fd_sc_hd__xnor2_1
XFILLER_67_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6813_ _6814_/A _6814_/B _6814_/C vssd1 vssd1 vccd1 vccd1 _6840_/A sky130_fd_sc_hd__a21oi_1
XFILLER_35_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3956_ _7223_/Q vssd1 vssd1 vccd1 vccd1 _5016_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6744_ _6744_/A _6744_/B vssd1 vssd1 vccd1 vccd1 _6782_/B sky130_fd_sc_hd__xor2_1
X_6675_ _6675_/A _6675_/B vssd1 vssd1 vccd1 vccd1 _6685_/A sky130_fd_sc_hd__nand2_1
X_3887_ _3887_/A _3887_/B vssd1 vssd1 vccd1 vccd1 _3889_/C sky130_fd_sc_hd__xnor2_1
X_5626_ _6624_/A _5985_/B vssd1 vssd1 vccd1 vccd1 _5627_/B sky130_fd_sc_hd__or2_1
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5557_ _5557_/A _5557_/B vssd1 vssd1 vccd1 vccd1 _5559_/A sky130_fd_sc_hd__or2_1
X_4508_ _4609_/A _4609_/B vssd1 vssd1 vccd1 vccd1 _4508_/Y sky130_fd_sc_hd__nand2_1
X_5488_ _6264_/A _5542_/B _5540_/A vssd1 vssd1 vccd1 vccd1 _5490_/C sky130_fd_sc_hd__mux2_1
X_4439_ _4439_/A _4439_/B vssd1 vssd1 vccd1 vccd1 _4440_/B sky130_fd_sc_hd__xor2_1
XFILLER_76_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7158_ _7225_/CLK _7158_/D vssd1 vssd1 vccd1 vccd1 _7158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7089_ _7089_/A _7093_/B vssd1 vssd1 vccd1 vccd1 _7089_/Y sky130_fd_sc_hd__nand2_1
X_6109_ _6109_/A _6110_/A vssd1 vssd1 vccd1 vccd1 _6111_/A sky130_fd_sc_hd__or2b_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4790_ _4790_/A _4790_/B vssd1 vssd1 vccd1 vccd1 _4791_/B sky130_fd_sc_hd__and2_1
XFILLER_60_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3810_ _3802_/Y _4485_/A _4633_/A vssd1 vssd1 vccd1 vccd1 _4339_/B sky130_fd_sc_hd__a21oi_1
XFILLER_20_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_29 _3672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3741_ _3742_/A vssd1 vssd1 vccd1 vccd1 _3741_/Y sky130_fd_sc_hd__inv_2
XANTENNA_18 _6194_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6460_ _6460_/A _6461_/A vssd1 vssd1 vccd1 vccd1 _6730_/A sky130_fd_sc_hd__or2b_1
XFILLER_9_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3672_ _3672_/A vssd1 vssd1 vccd1 vccd1 _3672_/Y sky130_fd_sc_hd__inv_2
X_6391_ _6391_/A hold6/X vssd1 vssd1 vccd1 vccd1 _6391_/X sky130_fd_sc_hd__or2_1
X_5411_ _5412_/B _5412_/C _6209_/A vssd1 vssd1 vccd1 vccd1 _5413_/A sky130_fd_sc_hd__a21oi_1
XFILLER_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5342_ _5339_/A _5218_/B _5341_/X vssd1 vssd1 vccd1 vccd1 _5381_/B sky130_fd_sc_hd__o21ba_1
XFILLER_101_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5273_ _5273_/A vssd1 vssd1 vccd1 vccd1 _7055_/A sky130_fd_sc_hd__clkbuf_2
X_7012_ _6990_/A _7005_/X _7011_/X _7007_/X vssd1 vssd1 vccd1 vccd1 _7183_/D sky130_fd_sc_hd__o211a_1
XFILLER_101_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4224_ _5019_/A _4328_/A _4225_/A _4326_/B vssd1 vssd1 vccd1 vccd1 _6722_/A sky130_fd_sc_hd__o22a_4
XFILLER_101_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4155_ _5017_/A _5017_/B vssd1 vssd1 vccd1 vccd1 _4157_/C sky130_fd_sc_hd__xnor2_1
XFILLER_55_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4086_ _7161_/Q vssd1 vssd1 vccd1 vccd1 _4572_/A sky130_fd_sc_hd__buf_2
XFILLER_36_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4988_ _5275_/A _5274_/A _7085_/A vssd1 vssd1 vccd1 vccd1 _4989_/B sky130_fd_sc_hd__and3_1
XFILLER_11_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3939_ _4412_/B vssd1 vssd1 vccd1 vccd1 _4799_/A sky130_fd_sc_hd__buf_2
X_6727_ _6727_/A _6727_/B _6457_/B vssd1 vssd1 vccd1 vccd1 _6767_/A sky130_fd_sc_hd__or3b_1
X_6658_ _6973_/A _6658_/B vssd1 vssd1 vccd1 vccd1 _6662_/A sky130_fd_sc_hd__xnor2_1
XFILLER_11_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5609_ _6564_/A vssd1 vssd1 vccd1 vccd1 _6571_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6589_ _6589_/A _6589_/B vssd1 vssd1 vccd1 vccd1 _6621_/B sky130_fd_sc_hd__xnor2_1
XFILLER_87_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput16 io_in[24] vssd1 vssd1 vccd1 vccd1 _6886_/C sky130_fd_sc_hd__buf_2
XFILLER_10_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7249__42 vssd1 vssd1 vccd1 vccd1 _7249__42/HI _7348_/A sky130_fd_sc_hd__conb_1
XFILLER_65_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5960_ _6665_/A vssd1 vssd1 vccd1 vccd1 _6693_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4911_ _4895_/A _4895_/C _4895_/D _4895_/B vssd1 vssd1 vccd1 vccd1 _4911_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5891_ _5894_/A _5894_/B _5890_/Y vssd1 vssd1 vccd1 vccd1 _6097_/B sky130_fd_sc_hd__a21oi_2
XFILLER_33_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4842_ _5644_/A _6678_/A vssd1 vssd1 vccd1 vccd1 _4910_/A sky130_fd_sc_hd__nand2_1
XFILLER_20_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4773_ _4816_/A _4816_/B vssd1 vssd1 vccd1 vccd1 _4817_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3724_ _3727_/A vssd1 vssd1 vccd1 vccd1 _3724_/Y sky130_fd_sc_hd__inv_2
X_6512_ _6541_/A _6510_/X _6541_/B vssd1 vssd1 vccd1 vccd1 _6512_/X sky130_fd_sc_hd__o21ba_1
X_6443_ _6443_/A _6491_/A vssd1 vssd1 vccd1 vccd1 _6443_/Y sky130_fd_sc_hd__nor2_1
X_3655_ _3679_/A vssd1 vssd1 vccd1 vccd1 _3660_/A sky130_fd_sc_hd__buf_8
XFILLER_9_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6374_ _6374_/A _6374_/B vssd1 vssd1 vccd1 vccd1 _6378_/A sky130_fd_sc_hd__xnor2_1
X_5325_ _5325_/A _5325_/B _5325_/C vssd1 vssd1 vccd1 vccd1 _5325_/X sky130_fd_sc_hd__and3_1
XFILLER_87_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5256_ _5256_/A _5263_/A vssd1 vssd1 vccd1 vccd1 _5257_/C sky130_fd_sc_hd__xnor2_1
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4207_ _6493_/C vssd1 vssd1 vccd1 vccd1 _6479_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_75_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5187_ _5037_/A _5037_/B _5036_/A vssd1 vssd1 vccd1 vccd1 _5364_/B sky130_fd_sc_hd__a21o_1
XFILLER_83_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4138_ _6794_/B _4138_/B vssd1 vssd1 vccd1 vccd1 _6617_/A sky130_fd_sc_hd__or2_2
X_4069_ _6445_/B _7160_/Q vssd1 vssd1 vccd1 vccd1 _4070_/B sky130_fd_sc_hd__and2b_1
XFILLER_73_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5110_ _5110_/A _5116_/B vssd1 vssd1 vccd1 vccd1 _5111_/C sky130_fd_sc_hd__xor2_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6090_ _6090_/A _6186_/A vssd1 vssd1 vccd1 vccd1 _6091_/B sky130_fd_sc_hd__xnor2_4
XFILLER_69_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _5243_/A _5041_/B vssd1 vssd1 vccd1 vccd1 _5096_/A sky130_fd_sc_hd__xnor2_2
XFILLER_97_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
X_6992_ _7052_/A vssd1 vssd1 vccd1 vccd1 _7045_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5943_ _5943_/A _5943_/B vssd1 vssd1 vccd1 vccd1 _5963_/A sky130_fd_sc_hd__or2_1
XFILLER_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5874_ _7014_/A _6480_/B vssd1 vssd1 vccd1 vccd1 _5912_/A sky130_fd_sc_hd__nand2_1
XFILLER_21_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4825_ _4870_/A _4870_/B _4824_/Y vssd1 vssd1 vccd1 vccd1 _4827_/B sky130_fd_sc_hd__a21o_1
X_4756_ _4756_/A _4756_/B vssd1 vssd1 vccd1 vccd1 _4782_/A sky130_fd_sc_hd__xnor2_1
X_3707_ _3709_/A vssd1 vssd1 vccd1 vccd1 _3707_/Y sky130_fd_sc_hd__inv_2
X_4687_ _4689_/A _4689_/B _4686_/Y vssd1 vssd1 vccd1 vccd1 _4720_/A sky130_fd_sc_hd__o21ai_1
X_3638_ _3641_/A vssd1 vssd1 vccd1 vccd1 _3638_/Y sky130_fd_sc_hd__inv_2
X_6426_ _6975_/A _6552_/A vssd1 vssd1 vccd1 vccd1 _6720_/A sky130_fd_sc_hd__nor2_1
X_6357_ _6316_/A _6357_/B vssd1 vssd1 vccd1 vccd1 _6357_/X sky130_fd_sc_hd__and2b_1
X_5308_ _5308_/A _5308_/B vssd1 vssd1 vccd1 vccd1 _5314_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6288_ _6546_/A vssd1 vssd1 vccd1 vccd1 _6528_/B sky130_fd_sc_hd__buf_2
X_5239_ _5239_/A _5239_/B vssd1 vssd1 vccd1 vccd1 _5240_/B sky130_fd_sc_hd__xnor2_2
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_47_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4610_ _7041_/A _4638_/B vssd1 vssd1 vccd1 vccd1 _4611_/B sky130_fd_sc_hd__nor2_1
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5590_ _5590_/A _5590_/B vssd1 vssd1 vccd1 vccd1 _5590_/X sky130_fd_sc_hd__or2_1
X_4541_ _7085_/A _4541_/B vssd1 vssd1 vccd1 vccd1 _4542_/B sky130_fd_sc_hd__nand2_1
X_4472_ _4472_/A _4472_/B vssd1 vssd1 vccd1 vccd1 _4564_/C sky130_fd_sc_hd__xnor2_1
X_7191_ _7222_/CLK _7191_/D vssd1 vssd1 vccd1 vccd1 _7191_/Q sky130_fd_sc_hd__dfxtp_1
X_6211_ _5450_/B _6127_/B _6210_/X vssd1 vssd1 vccd1 vccd1 _6262_/B sky130_fd_sc_hd__a21o_1
X_6142_ _7009_/A _6142_/B vssd1 vssd1 vccd1 vccd1 _6142_/X sky130_fd_sc_hd__and2b_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6073_ _6073_/A _6073_/B vssd1 vssd1 vccd1 vccd1 _6167_/B sky130_fd_sc_hd__nand2_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _5022_/Y _5171_/A vssd1 vssd1 vccd1 vccd1 _5024_/X sky130_fd_sc_hd__and2b_1
XFILLER_38_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6975_ _6975_/A _6975_/B vssd1 vssd1 vccd1 vccd1 _6975_/X sky130_fd_sc_hd__or2_1
XFILLER_53_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5926_ _5926_/A _5943_/A vssd1 vssd1 vccd1 vccd1 _5927_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5857_ _5857_/A _5857_/B vssd1 vssd1 vccd1 vccd1 _5859_/C sky130_fd_sc_hd__xnor2_1
X_4808_ _4808_/A _4808_/B vssd1 vssd1 vccd1 vccd1 _4810_/A sky130_fd_sc_hd__xnor2_1
XFILLER_21_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5788_ _6070_/A _5788_/B vssd1 vssd1 vccd1 vccd1 _6065_/A sky130_fd_sc_hd__nand2_1
X_4739_ _4739_/A _4739_/B vssd1 vssd1 vccd1 vccd1 _4754_/B sky130_fd_sc_hd__xor2_1
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6409_ _6409_/A _6409_/B vssd1 vssd1 vccd1 vccd1 _6559_/A sky130_fd_sc_hd__xnor2_1
X_7389_ _7389_/A _3681_/Y vssd1 vssd1 vccd1 vccd1 io_out[31] sky130_fd_sc_hd__ebufn_8
X_7303__96 vssd1 vssd1 vccd1 vccd1 _7303__96/HI _7411_/A sky130_fd_sc_hd__conb_1
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6760_ _6812_/A _6760_/B vssd1 vssd1 vccd1 vccd1 _6777_/A sky130_fd_sc_hd__nor2_1
XFILLER_23_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5711_ hold89/A _5749_/A vssd1 vssd1 vccd1 vccd1 _5714_/A sky130_fd_sc_hd__nand2_2
X_3972_ _5023_/A _3972_/B vssd1 vssd1 vccd1 vccd1 _3974_/B sky130_fd_sc_hd__or2_1
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6691_ _6691_/A _6691_/B vssd1 vssd1 vccd1 vccd1 _6691_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5642_ _6794_/A _6087_/B vssd1 vssd1 vccd1 vccd1 _5643_/A sky130_fd_sc_hd__nand2_1
X_5573_ hold14/X vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__inv_2
X_4524_ _4444_/A _4444_/B _4523_/Y vssd1 vssd1 vccd1 vccd1 _5104_/A sky130_fd_sc_hd__a21oi_1
X_4455_ _4453_/A _4666_/A _4556_/A vssd1 vssd1 vccd1 vccd1 _4472_/A sky130_fd_sc_hd__a21oi_1
X_4386_ _4304_/A _4304_/B _4385_/X vssd1 vssd1 vccd1 vccd1 _5043_/B sky130_fd_sc_hd__a21oi_2
X_7174_ _7183_/CLK _7174_/D vssd1 vssd1 vccd1 vccd1 _7174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6125_ _6125_/A _6125_/B vssd1 vssd1 vccd1 vccd1 _6210_/B sky130_fd_sc_hd__nor2_2
XFILLER_100_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ _6057_/A _6057_/B vssd1 vssd1 vccd1 vccd1 _6056_/Y sky130_fd_sc_hd__nand2_1
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5007_ _4143_/X _5004_/Y _5006_/Y vssd1 vssd1 vccd1 vccd1 _5015_/A sky130_fd_sc_hd__o21ai_2
XFILLER_81_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6958_ _7095_/A vssd1 vssd1 vccd1 vccd1 _7114_/B sky130_fd_sc_hd__clkbuf_2
X_5909_ _5824_/A _5749_/A _5880_/C vssd1 vssd1 vccd1 vccd1 _5910_/B sky130_fd_sc_hd__o21ba_1
X_6889_ _6889_/A vssd1 vssd1 vccd1 vccd1 _6893_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4240_ _4240_/A _4240_/B _4240_/C vssd1 vssd1 vccd1 vccd1 _4260_/A sky130_fd_sc_hd__and3_1
XFILLER_101_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4171_ _4873_/A _3922_/B _3873_/A vssd1 vssd1 vccd1 vccd1 _4174_/B sky130_fd_sc_hd__a21bo_1
XFILLER_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7294__87 vssd1 vssd1 vccd1 vccd1 _7294__87/HI _7402_/A sky130_fd_sc_hd__conb_1
XFILLER_82_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6812_ _6812_/A _6812_/B vssd1 vssd1 vccd1 vccd1 _6814_/C sky130_fd_sc_hd__xnor2_1
XFILLER_35_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3955_ _6484_/A _7223_/Q vssd1 vssd1 vccd1 vccd1 _4154_/A sky130_fd_sc_hd__nand2b_2
X_6743_ _6743_/A _6743_/B vssd1 vssd1 vccd1 vccd1 _6744_/B sky130_fd_sc_hd__nand2_1
X_6674_ _6674_/A _6674_/B vssd1 vssd1 vccd1 vccd1 _6675_/B sky130_fd_sc_hd__or2_1
XFILLER_31_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3886_ _3886_/A _3886_/B vssd1 vssd1 vccd1 vccd1 _3887_/B sky130_fd_sc_hd__nor2_1
X_5625_ _5625_/A _5625_/B vssd1 vssd1 vccd1 vccd1 _5736_/C sky130_fd_sc_hd__nand2_1
X_5556_ _5556_/A _5556_/B _5556_/C vssd1 vssd1 vccd1 vccd1 _5557_/B sky130_fd_sc_hd__nor3_1
X_4507_ _4507_/A _4507_/B vssd1 vssd1 vccd1 vccd1 _4609_/B sky130_fd_sc_hd__xnor2_1
X_5487_ _6966_/A _5143_/X _5486_/Y vssd1 vssd1 vccd1 vccd1 _5540_/A sky130_fd_sc_hd__a21o_1
X_4438_ _4548_/A _4548_/B _4437_/X vssd1 vssd1 vccd1 vccd1 _4492_/B sky130_fd_sc_hd__o21a_1
X_7226_ _7226_/CLK _7226_/D vssd1 vssd1 vccd1 vccd1 _7391_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_98_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7157_ _7172_/CLK _7157_/D vssd1 vssd1 vccd1 vccd1 _7157_/Q sky130_fd_sc_hd__dfxtp_1
X_4369_ _4949_/A _4369_/B vssd1 vssd1 vccd1 vccd1 _4388_/A sky130_fd_sc_hd__xor2_4
XFILLER_100_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7088_ _7101_/A vssd1 vssd1 vccd1 vccd1 _7088_/X sky130_fd_sc_hd__clkbuf_2
X_6108_ _6108_/A _6108_/B vssd1 vssd1 vccd1 vccd1 _6115_/A sky130_fd_sc_hd__nand2_2
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6039_ _5688_/B _6039_/B _6045_/B vssd1 vssd1 vccd1 vccd1 _6039_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_39_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_19 _6943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3740_ _3742_/A vssd1 vssd1 vccd1 vccd1 _3740_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3671_ _3672_/A vssd1 vssd1 vccd1 vccd1 _3671_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6390_ _6390_/A _6390_/B vssd1 vssd1 vccd1 vccd1 _6390_/X sky130_fd_sc_hd__xor2_1
X_5410_ _6129_/A vssd1 vssd1 vccd1 vccd1 _6209_/A sky130_fd_sc_hd__clkbuf_2
X_5341_ _5341_/A _5341_/B _5341_/C vssd1 vssd1 vccd1 vccd1 _5341_/X sky130_fd_sc_hd__and3_1
X_7011_ _7011_/A _7011_/B vssd1 vssd1 vccd1 vccd1 _7011_/X sky130_fd_sc_hd__or2_1
X_5272_ _5386_/B _5271_/Y vssd1 vssd1 vccd1 vccd1 _5282_/A sky130_fd_sc_hd__or2b_1
X_4223_ _4794_/A _5972_/C _6719_/B vssd1 vssd1 vccd1 vccd1 _4326_/B sky130_fd_sc_hd__a21oi_4
XFILLER_101_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4154_ _4154_/A _4154_/B vssd1 vssd1 vccd1 vccd1 _5017_/B sky130_fd_sc_hd__xnor2_1
XFILLER_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4085_ _7166_/Q vssd1 vssd1 vccd1 vccd1 _5002_/A sky130_fd_sc_hd__buf_2
XFILLER_36_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6726_ _6765_/B _6726_/B vssd1 vssd1 vccd1 vccd1 _6727_/B sky130_fd_sc_hd__nand2_1
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4987_ _4987_/A vssd1 vssd1 vccd1 vccd1 _4989_/A sky130_fd_sc_hd__inv_2
X_3938_ _5274_/A _3995_/A vssd1 vssd1 vccd1 vccd1 _3942_/A sky130_fd_sc_hd__nor2_1
X_3869_ _7210_/Q vssd1 vssd1 vccd1 vccd1 _7083_/A sky130_fd_sc_hd__inv_2
X_6657_ _6657_/A _6624_/X vssd1 vssd1 vccd1 vccd1 _6658_/B sky130_fd_sc_hd__or2b_1
X_6588_ _6588_/A _6588_/B vssd1 vssd1 vccd1 vccd1 _6589_/B sky130_fd_sc_hd__xnor2_4
XFILLER_11_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5608_ _6067_/A vssd1 vssd1 vccd1 vccd1 _5801_/A sky130_fd_sc_hd__buf_2
XFILLER_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5539_ _5479_/A _5479_/B _5538_/X vssd1 vssd1 vccd1 vccd1 _5584_/A sky130_fd_sc_hd__o21bai_2
XFILLER_87_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7209_ _7221_/CLK _7209_/D vssd1 vssd1 vccd1 vccd1 _7209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput17 io_in[8] vssd1 vssd1 vccd1 vccd1 _7117_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_6_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7264__57 vssd1 vssd1 vccd1 vccd1 _7264__57/HI _7363_/A sky130_fd_sc_hd__conb_1
XFILLER_92_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4910_ _4910_/A _4910_/B vssd1 vssd1 vccd1 vccd1 _4910_/X sky130_fd_sc_hd__and2_1
XFILLER_73_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5890_ _5890_/A _5890_/B vssd1 vssd1 vccd1 vccd1 _5890_/Y sky130_fd_sc_hd__nor2_1
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4841_ _6480_/B vssd1 vssd1 vccd1 vccd1 _6678_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4772_ _4772_/A _4772_/B vssd1 vssd1 vccd1 vccd1 _4816_/B sky130_fd_sc_hd__xnor2_1
XFILLER_20_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6511_ _6506_/A _6506_/B _6506_/C vssd1 vssd1 vccd1 vccd1 _6541_/B sky130_fd_sc_hd__a21oi_1
X_3723_ _3727_/A vssd1 vssd1 vccd1 vccd1 _3723_/Y sky130_fd_sc_hd__inv_2
X_6442_ _6443_/A _6491_/A vssd1 vssd1 vccd1 vccd1 _6481_/B sky130_fd_sc_hd__xor2_2
XFILLER_9_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3654_ input1/X vssd1 vssd1 vccd1 vccd1 _3679_/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_3_0_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7224_/CLK
+ sky130_fd_sc_hd__clkbuf_2
X_6373_ _6341_/A _6341_/B _6372_/X vssd1 vssd1 vccd1 vccd1 _6374_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5324_ _5239_/A _5239_/B _5323_/X vssd1 vssd1 vccd1 vccd1 _5359_/A sky130_fd_sc_hd__a21bo_1
X_5255_ _5107_/A _5107_/B _5254_/X vssd1 vssd1 vccd1 vccd1 _5263_/A sky130_fd_sc_hd__o21ba_1
X_4206_ _7153_/Q vssd1 vssd1 vccd1 vccd1 _6493_/C sky130_fd_sc_hd__inv_2
XFILLER_68_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5186_ _5093_/A _5093_/B _5092_/A vssd1 vssd1 vccd1 vccd1 _5365_/B sky130_fd_sc_hd__a21o_2
XFILLER_95_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4137_ _5002_/A _4279_/A _5167_/A vssd1 vssd1 vccd1 vccd1 _6794_/B sky130_fd_sc_hd__and3_1
X_4068_ hold94/A _6507_/A vssd1 vssd1 vccd1 vccd1 _4215_/A sky130_fd_sc_hd__and2_1
XFILLER_43_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6709_ _6261_/X _6707_/X hold50/X _6196_/X vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__o211a_1
XFILLER_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _4167_/A _4167_/B _5039_/X vssd1 vssd1 vccd1 vccd1 _5041_/B sky130_fd_sc_hd__a21bo_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6991_ _6969_/A _6977_/X _6990_/X _6979_/X vssd1 vssd1 vccd1 vccd1 _7175_/D sky130_fd_sc_hd__o211a_1
X_5942_ _5942_/A _5942_/B vssd1 vssd1 vccd1 vccd1 _5943_/B sky130_fd_sc_hd__and2_1
XFILLER_53_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5873_ _5873_/A _6480_/B vssd1 vssd1 vccd1 vccd1 _5912_/B sky130_fd_sc_hd__or2_1
X_4824_ _4824_/A _4872_/A vssd1 vssd1 vccd1 vccd1 _4824_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4755_ _4757_/A _4757_/B _4754_/Y vssd1 vssd1 vccd1 vccd1 _4788_/A sky130_fd_sc_hd__o21ai_1
XFILLER_21_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3706_ _3709_/A vssd1 vssd1 vccd1 vccd1 _3706_/Y sky130_fd_sc_hd__inv_2
X_4686_ _4686_/A _4686_/B vssd1 vssd1 vccd1 vccd1 _4686_/Y sky130_fd_sc_hd__nand2_1
X_6425_ _6528_/A _6528_/B vssd1 vssd1 vccd1 vccd1 _6552_/A sky130_fd_sc_hd__nand2_1
X_3637_ _3641_/A vssd1 vssd1 vccd1 vccd1 _3637_/Y sky130_fd_sc_hd__inv_2
X_6356_ _6356_/A _6388_/B vssd1 vssd1 vccd1 vccd1 _6359_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5307_ _5307_/A _5307_/B vssd1 vssd1 vccd1 vccd1 _5308_/B sky130_fd_sc_hd__and2_1
X_6287_ _5801_/A _6289_/B _6230_/B vssd1 vssd1 vccd1 vccd1 _6294_/B sky130_fd_sc_hd__o21bai_1
XFILLER_76_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5238_ _5238_/A _5323_/A vssd1 vssd1 vccd1 vccd1 _5239_/B sky130_fd_sc_hd__xnor2_1
XFILLER_68_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5169_ _5167_/A _6464_/A _5168_/A vssd1 vssd1 vccd1 vccd1 _5169_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_68_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7313__106 vssd1 vssd1 vccd1 vccd1 _7313__106/HI _7421_/A sky130_fd_sc_hd__conb_1
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_7234__27 vssd1 vssd1 vccd1 vccd1 _7234__27/HI _7333_/A sky130_fd_sc_hd__conb_1
XFILLER_47_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4540_ _4649_/A _4540_/B _4541_/B vssd1 vssd1 vccd1 vccd1 _4542_/A sky130_fd_sc_hd__or3_1
X_4471_ _4569_/A _4569_/B vssd1 vssd1 vccd1 vccd1 _4564_/B sky130_fd_sc_hd__and2b_1
XFILLER_7_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7190_ _7222_/CLK _7190_/D vssd1 vssd1 vccd1 vccd1 _7190_/Q sky130_fd_sc_hd__dfxtp_1
X_6210_ _6210_/A _6210_/B vssd1 vssd1 vccd1 vccd1 _6210_/X sky130_fd_sc_hd__and2_1
X_6141_ _6142_/B _7009_/A vssd1 vssd1 vccd1 vccd1 _6141_/X sky130_fd_sc_hd__and2b_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6072_ _6073_/A _6073_/B vssd1 vssd1 vccd1 vccd1 _6074_/A sky130_fd_sc_hd__or2_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5023_ _5023_/A _5023_/B vssd1 vssd1 vccd1 vccd1 _5171_/A sky130_fd_sc_hd__nand2_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6974_ _6950_/A _6964_/X _6973_/Y _6967_/X vssd1 vssd1 vccd1 vccd1 _7169_/D sky130_fd_sc_hd__o211a_1
XFILLER_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5925_ _5942_/A _5942_/B vssd1 vssd1 vccd1 vccd1 _5943_/A sky130_fd_sc_hd__nor2_1
XFILLER_41_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5856_ _5856_/A _5856_/B vssd1 vssd1 vccd1 vccd1 _5857_/B sky130_fd_sc_hd__nor2_1
X_4807_ _4815_/A _4815_/B _4806_/A vssd1 vssd1 vccd1 vccd1 _4809_/A sky130_fd_sc_hd__a21o_1
XFILLER_21_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5787_ _5787_/A _5787_/B _5787_/C vssd1 vssd1 vccd1 vccd1 _5788_/B sky130_fd_sc_hd__nand3_1
X_4738_ _4759_/A _4759_/B _4737_/A vssd1 vssd1 vccd1 vccd1 _4754_/A sky130_fd_sc_hd__o21ai_1
X_4669_ _4723_/A _4723_/B vssd1 vssd1 vccd1 vccd1 _4676_/A sky130_fd_sc_hd__and2_1
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6408_ _6613_/A _6613_/B _6704_/B vssd1 vssd1 vccd1 vccd1 _6586_/B sky130_fd_sc_hd__a21oi_2
X_7388_ _7388_/A _3680_/Y vssd1 vssd1 vccd1 vccd1 io_out[30] sky130_fd_sc_hd__ebufn_8
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6339_ _6413_/A _6420_/B vssd1 vssd1 vccd1 vccd1 _6375_/B sky130_fd_sc_hd__nand2_1
XFILLER_95_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3971_ _5016_/A _6022_/A vssd1 vssd1 vccd1 vccd1 _3972_/B sky130_fd_sc_hd__and2b_1
X_5710_ _5710_/A _5710_/B vssd1 vssd1 vccd1 vccd1 _6057_/A sky130_fd_sc_hd__xnor2_4
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6690_ _6690_/A _6690_/B vssd1 vssd1 vccd1 vccd1 _6691_/B sky130_fd_sc_hd__xnor2_1
X_5641_ _6061_/B vssd1 vssd1 vccd1 vccd1 _6794_/A sky130_fd_sc_hd__buf_2
XFILLER_31_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5572_ _5262_/X _5570_/Y hold60/X _7226_/D vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__o211a_1
X_4523_ _4523_/A _4523_/B vssd1 vssd1 vccd1 vccd1 _4523_/Y sky130_fd_sc_hd__nor2_1
X_4454_ _4555_/A _4555_/B vssd1 vssd1 vccd1 vccd1 _4556_/A sky130_fd_sc_hd__nor2_1
X_4385_ _4303_/A _4385_/B vssd1 vssd1 vccd1 vccd1 _4385_/X sky130_fd_sc_hd__and2b_1
X_7173_ _7183_/CLK _7173_/D vssd1 vssd1 vccd1 vccd1 _7173_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6124_ _6124_/A _6124_/B _6124_/C vssd1 vssd1 vccd1 vccd1 _6125_/B sky130_fd_sc_hd__nor3_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _6055_/A _6055_/B vssd1 vssd1 vccd1 vccd1 _6171_/A sky130_fd_sc_hd__xnor2_2
XFILLER_85_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5006_ _5406_/A _5006_/B vssd1 vssd1 vccd1 vccd1 _5006_/Y sky130_fd_sc_hd__nand2_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6957_ _6588_/A _6949_/X _6956_/Y _6952_/X vssd1 vssd1 vccd1 vccd1 _7163_/D sky130_fd_sc_hd__o211a_1
XFILLER_53_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5908_ _5908_/A _5908_/B vssd1 vssd1 vccd1 vccd1 _5924_/A sky130_fd_sc_hd__xnor2_1
X_6888_ _6891_/B _6891_/C input9/X vssd1 vssd1 vccd1 vccd1 _6889_/A sky130_fd_sc_hd__and3b_1
X_5839_ _5839_/A _5839_/B vssd1 vssd1 vccd1 vccd1 _5868_/A sky130_fd_sc_hd__or2_1
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7319__112 vssd1 vssd1 vccd1 vccd1 _7319__112/HI _7427_/A sky130_fd_sc_hd__conb_1
XFILLER_29_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4170_ _4392_/B vssd1 vssd1 vccd1 vccd1 _7043_/A sky130_fd_sc_hd__buf_2
XFILLER_82_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6811_ _6837_/A _6837_/B vssd1 vssd1 vccd1 vccd1 _6812_/B sky130_fd_sc_hd__xor2_1
X_3954_ _7157_/Q vssd1 vssd1 vccd1 vccd1 _6484_/A sky130_fd_sc_hd__clkbuf_2
X_6742_ _6778_/A _6778_/B _6778_/C vssd1 vssd1 vccd1 vccd1 _6743_/B sky130_fd_sc_hd__or3_1
X_3885_ _5129_/A _3910_/A _4957_/A vssd1 vssd1 vccd1 vccd1 _3886_/B sky130_fd_sc_hd__a21oi_1
XFILLER_31_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6673_ _6960_/A _6704_/B _6704_/C vssd1 vssd1 vccd1 vccd1 _6673_/X sky130_fd_sc_hd__a21o_1
X_5624_ _5736_/B vssd1 vssd1 vccd1 vccd1 _6659_/A sky130_fd_sc_hd__buf_2
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5555_ _5556_/A _5556_/B _5556_/C vssd1 vssd1 vccd1 vccd1 _5557_/A sky130_fd_sc_hd__o21a_1
X_4506_ _4506_/A _4506_/B _4506_/C vssd1 vssd1 vccd1 vccd1 _4507_/B sky130_fd_sc_hd__and3_1
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5486_ _6524_/A _5486_/B vssd1 vssd1 vccd1 vccd1 _5486_/Y sky130_fd_sc_hd__nand2_1
X_4437_ _4437_/A _4437_/B vssd1 vssd1 vccd1 vccd1 _4437_/X sky130_fd_sc_hd__or2_1
X_7225_ _7225_/CLK _7225_/D vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__dfxtp_1
X_7156_ _7225_/CLK _7156_/D vssd1 vssd1 vccd1 vccd1 _7156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6107_ _6107_/A _6107_/B vssd1 vssd1 vccd1 vccd1 _6108_/B sky130_fd_sc_hd__or2_1
XFILLER_58_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4368_ _4285_/A _3797_/B _4367_/X vssd1 vssd1 vccd1 vccd1 _4369_/B sky130_fd_sc_hd__a21bo_1
X_7087_ hold58/X _7075_/X _7085_/Y _7086_/X vssd1 vssd1 vccd1 vccd1 _7211_/D sky130_fd_sc_hd__o211a_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4299_ _4374_/A _4124_/A _4298_/Y vssd1 vssd1 vccd1 vccd1 _4300_/B sky130_fd_sc_hd__o21a_1
X_6038_ _6132_/A _6038_/B vssd1 vssd1 vccd1 vccd1 _6147_/B sky130_fd_sc_hd__xnor2_4
XFILLER_39_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3670_ _3672_/A vssd1 vssd1 vccd1 vccd1 _3670_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5340_ _5340_/A _5446_/C vssd1 vssd1 vccd1 vccd1 _5381_/A sky130_fd_sc_hd__xor2_1
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5271_ _5271_/A _5271_/B vssd1 vssd1 vccd1 vccd1 _5271_/Y sky130_fd_sc_hd__nand2_1
X_4222_ _4795_/A _7163_/Q vssd1 vssd1 vccd1 vccd1 _6719_/B sky130_fd_sc_hd__and2b_2
X_7010_ _6852_/A _7005_/X _7009_/X _7007_/X vssd1 vssd1 vccd1 vccd1 _7182_/D sky130_fd_sc_hd__o211a_1
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4153_ _5019_/A _6016_/A vssd1 vssd1 vccd1 vccd1 _4154_/B sky130_fd_sc_hd__xnor2_1
X_4084_ _4084_/A _4084_/B vssd1 vssd1 vccd1 vccd1 _4202_/A sky130_fd_sc_hd__nor2_2
XFILLER_36_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4986_ _5275_/A _4986_/B vssd1 vssd1 vccd1 vccd1 _4987_/A sky130_fd_sc_hd__or2_1
XFILLER_23_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3937_ _5274_/A _3944_/B _3936_/X vssd1 vssd1 vccd1 vccd1 _4026_/A sky130_fd_sc_hd__a21o_2
X_6725_ _6725_/A _6725_/B vssd1 vssd1 vccd1 vccd1 _6726_/B sky130_fd_sc_hd__or2_1
XFILLER_51_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3868_ _7213_/Q vssd1 vssd1 vccd1 vccd1 _5131_/A sky130_fd_sc_hd__clkbuf_2
X_6656_ _6656_/A _6656_/B vssd1 vssd1 vccd1 vccd1 _6664_/A sky130_fd_sc_hd__or2_1
X_6587_ _6931_/A _6479_/B _6678_/A vssd1 vssd1 vccd1 vccd1 _6588_/B sky130_fd_sc_hd__a21oi_2
X_3799_ _4339_/A vssd1 vssd1 vccd1 vccd1 _3811_/A sky130_fd_sc_hd__inv_2
X_5607_ _5802_/A _5607_/B vssd1 vssd1 vccd1 vccd1 _5801_/B sky130_fd_sc_hd__or2_2
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5538_ _5493_/A _5538_/B vssd1 vssd1 vccd1 vccd1 _5538_/X sky130_fd_sc_hd__and2b_1
X_7208_ _7221_/CLK _7208_/D vssd1 vssd1 vccd1 vccd1 _7208_/Q sky130_fd_sc_hd__dfxtp_1
X_5469_ _5371_/A _5371_/B _5468_/X vssd1 vssd1 vccd1 vccd1 _5475_/B sky130_fd_sc_hd__o21ai_2
XFILLER_59_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7139_ _7151_/CLK hold36/X vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__dfxtp_1
XFILLER_86_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 io_in[9] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4840_ _5691_/B vssd1 vssd1 vccd1 vccd1 _6480_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4771_ _4771_/A _4771_/B vssd1 vssd1 vccd1 vccd1 _4816_/A sky130_fd_sc_hd__or2_1
X_6510_ _6506_/C _6565_/A _6542_/B vssd1 vssd1 vccd1 vccd1 _6510_/X sky130_fd_sc_hd__and3b_1
X_3722_ _3734_/A vssd1 vssd1 vccd1 vccd1 _3727_/A sky130_fd_sc_hd__buf_12
XFILLER_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6441_ _6441_/A _6441_/B _6441_/C _6441_/D vssd1 vssd1 vccd1 vccd1 _6491_/A sky130_fd_sc_hd__or4_2
X_3653_ _3653_/A vssd1 vssd1 vccd1 vccd1 _3653_/Y sky130_fd_sc_hd__inv_2
X_6372_ _6338_/B _6372_/B vssd1 vssd1 vccd1 vccd1 _6372_/X sky130_fd_sc_hd__and2b_1
X_5323_ _5323_/A _5238_/A vssd1 vssd1 vccd1 vccd1 _5323_/X sky130_fd_sc_hd__or2b_1
XFILLER_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5254_ _5106_/A _5254_/B vssd1 vssd1 vccd1 vccd1 _5254_/X sky130_fd_sc_hd__and2b_1
X_4205_ _6110_/A vssd1 vssd1 vccd1 vccd1 _4429_/A sky130_fd_sc_hd__clkbuf_4
X_5185_ _5361_/A _5361_/B vssd1 vssd1 vccd1 vccd1 _5242_/A sky130_fd_sc_hd__xnor2_2
X_4136_ _5021_/A vssd1 vssd1 vccd1 vccd1 _5167_/A sky130_fd_sc_hd__buf_2
XFILLER_95_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4067_ _6494_/B vssd1 vssd1 vccd1 vccd1 _6507_/A sky130_fd_sc_hd__inv_2
XFILLER_24_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4969_ _5133_/A _5292_/A vssd1 vssd1 vccd1 vccd1 _5146_/B sky130_fd_sc_hd__and2_1
XFILLER_11_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6708_ _6845_/A hold51/X vssd1 vssd1 vccd1 vccd1 hold50/A sky130_fd_sc_hd__or2_1
X_6639_ _6639_/A _6639_/B vssd1 vssd1 vccd1 vccd1 _6641_/B sky130_fd_sc_hd__xor2_2
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6990_ _6990_/A _7011_/B vssd1 vssd1 vccd1 vccd1 _6990_/X sky130_fd_sc_hd__or2_1
XFILLER_92_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5941_ _5941_/A _5941_/B vssd1 vssd1 vccd1 vccd1 _5967_/A sky130_fd_sc_hd__xor2_1
XFILLER_25_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5872_ _5872_/A _5872_/B vssd1 vssd1 vccd1 vccd1 _5876_/A sky130_fd_sc_hd__xnor2_2
XFILLER_61_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4823_ _4824_/A _4872_/A vssd1 vssd1 vccd1 vccd1 _4870_/B sky130_fd_sc_hd__xor2_2
XFILLER_61_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4754_ _4754_/A _4754_/B vssd1 vssd1 vccd1 vccd1 _4754_/Y sky130_fd_sc_hd__nand2_1
X_3705_ _3709_/A vssd1 vssd1 vccd1 vccd1 _3705_/Y sky130_fd_sc_hd__inv_2
X_4685_ _4739_/A _4739_/B _4684_/Y _4678_/B vssd1 vssd1 vccd1 vccd1 _4689_/B sky130_fd_sc_hd__o2bb2a_1
X_3636_ _3648_/A vssd1 vssd1 vccd1 vccd1 _3641_/A sky130_fd_sc_hd__buf_12
X_6424_ _6424_/A _6423_/Y vssd1 vssd1 vccd1 vccd1 _6718_/A sky130_fd_sc_hd__or2b_1
X_6355_ _6313_/A _6313_/B _6354_/X vssd1 vssd1 vccd1 vccd1 _6388_/B sky130_fd_sc_hd__a21bo_1
X_6286_ _6537_/B _6286_/B vssd1 vssd1 vccd1 vccd1 _6289_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5306_ _5307_/A _5307_/B vssd1 vssd1 vccd1 vccd1 _5308_/A sky130_fd_sc_hd__nor2_1
XFILLER_88_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5237_ _5088_/A _5088_/B _5236_/X vssd1 vssd1 vccd1 vccd1 _5323_/A sky130_fd_sc_hd__a21oi_2
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5168_ _5168_/A _6464_/A vssd1 vssd1 vccd1 vccd1 _5168_/X sky130_fd_sc_hd__or2_1
X_4119_ _4202_/A _4202_/B _4084_/A vssd1 vssd1 vccd1 vccd1 _4166_/A sky130_fd_sc_hd__a21o_2
X_5099_ _5097_/Y _4391_/B _5098_/Y vssd1 vssd1 vccd1 vccd1 _5100_/B sky130_fd_sc_hd__a21oi_4
XFILLER_29_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_47_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4470_ _4566_/A _4470_/B vssd1 vssd1 vccd1 vccd1 _4569_/B sky130_fd_sc_hd__xnor2_1
XFILLER_7_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6140_ _6140_/A vssd1 vssd1 vccd1 vccd1 _7009_/A sky130_fd_sc_hd__buf_2
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6071_ _6167_/A _6071_/B vssd1 vssd1 vccd1 vccd1 _6073_/B sky130_fd_sc_hd__and2_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5022_ _5023_/A _5023_/B vssd1 vssd1 vccd1 vccd1 _5022_/Y sky130_fd_sc_hd__nor2_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6973_ _6973_/A _6983_/B vssd1 vssd1 vccd1 vccd1 _6973_/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5924_ _5924_/A _5924_/B vssd1 vssd1 vccd1 vccd1 _5942_/B sky130_fd_sc_hd__xor2_1
XFILLER_34_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5855_ _6560_/A _5808_/B _5807_/B _6413_/B vssd1 vssd1 vccd1 vccd1 _5856_/B sky130_fd_sc_hd__o211a_1
X_4806_ _4806_/A _4806_/B vssd1 vssd1 vccd1 vccd1 _4815_/B sky130_fd_sc_hd__nor2_1
X_5786_ _5787_/A _5787_/B _5787_/C vssd1 vssd1 vccd1 vccd1 _6070_/A sky130_fd_sc_hd__a21o_1
X_4737_ _4737_/A _4737_/B vssd1 vssd1 vccd1 vccd1 _4759_/B sky130_fd_sc_hd__nand2_1
X_4668_ _4674_/A _4668_/B vssd1 vssd1 vccd1 vccd1 _4723_/B sky130_fd_sc_hd__xnor2_1
X_3619_ _3622_/A vssd1 vssd1 vccd1 vccd1 _3619_/Y sky130_fd_sc_hd__inv_2
X_6407_ _6956_/A _4330_/A _6698_/A vssd1 vssd1 vccd1 vccd1 _6613_/B sky130_fd_sc_hd__o21ai_2
X_4599_ _4599_/A _4599_/B vssd1 vssd1 vccd1 vccd1 _4629_/A sky130_fd_sc_hd__xnor2_1
X_7387_ _7387_/A _3678_/Y vssd1 vssd1 vccd1 vccd1 io_out[29] sky130_fd_sc_hd__ebufn_8
X_6338_ _6372_/B _6338_/B vssd1 vssd1 vccd1 vccd1 _6341_/A sky130_fd_sc_hd__xnor2_1
XFILLER_95_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6269_ _6269_/A _6854_/A vssd1 vssd1 vccd1 vccd1 _6270_/B sky130_fd_sc_hd__nand2_1
XFILLER_48_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3970_ _7158_/Q vssd1 vssd1 vccd1 vccd1 _6022_/A sky130_fd_sc_hd__buf_2
XFILLER_31_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5640_ _5640_/A vssd1 vssd1 vccd1 vccd1 _6061_/B sky130_fd_sc_hd__clkbuf_2
X_5571_ _5594_/A hold61/X vssd1 vssd1 vccd1 vccd1 hold60/A sky130_fd_sc_hd__or2_1
XFILLER_31_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4522_ _4522_/A _4522_/B vssd1 vssd1 vccd1 vccd1 _4525_/A sky130_fd_sc_hd__xor2_1
X_4453_ _4453_/A _4666_/A vssd1 vssd1 vccd1 vccd1 _4555_/B sky130_fd_sc_hd__xnor2_1
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7172_ _7172_/CLK _7172_/D vssd1 vssd1 vccd1 vccd1 _7172_/Q sky130_fd_sc_hd__dfxtp_1
X_4384_ _4384_/A _4384_/B vssd1 vssd1 vccd1 vccd1 _5043_/A sky130_fd_sc_hd__xnor2_2
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6123_ _6124_/A _6124_/C _6124_/B vssd1 vssd1 vccd1 vccd1 _6125_/A sky130_fd_sc_hd__o21a_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ _6054_/A _6054_/B vssd1 vssd1 vccd1 vccd1 _6055_/B sky130_fd_sc_hd__xnor2_2
XFILLER_39_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _5784_/B vssd1 vssd1 vccd1 vccd1 _5406_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_66_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6956_ _6956_/A _6956_/B vssd1 vssd1 vccd1 vccd1 _6956_/Y sky130_fd_sc_hd__nand2_1
XFILLER_26_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5907_ _5907_/A _5907_/B vssd1 vssd1 vccd1 vccd1 _5928_/B sky130_fd_sc_hd__xor2_1
XFILLER_53_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6887_ _6887_/A _6887_/B _6887_/C vssd1 vssd1 vccd1 vccd1 _6891_/C sky130_fd_sc_hd__nor3_1
X_5838_ _5813_/B _5838_/B vssd1 vssd1 vccd1 vccd1 _5839_/B sky130_fd_sc_hd__and2b_1
X_5769_ _5770_/A _5770_/B vssd1 vssd1 vccd1 vccd1 _5826_/B sky130_fd_sc_hd__xnor2_1
XFILLER_22_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6810_ _6777_/A _6777_/B _6809_/Y vssd1 vssd1 vccd1 vccd1 _6837_/B sky130_fd_sc_hd__a21bo_1
XFILLER_63_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3953_ hold94/A _4036_/A vssd1 vssd1 vccd1 vccd1 _4157_/A sky130_fd_sc_hd__or2_1
X_6741_ _6778_/A _6778_/B _6778_/C vssd1 vssd1 vccd1 vccd1 _6743_/A sky130_fd_sc_hd__o21ai_1
XFILLER_35_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6672_ _6672_/A _6672_/B vssd1 vssd1 vccd1 vccd1 _6704_/C sky130_fd_sc_hd__nor2_1
X_3884_ _5129_/A _3910_/A _4957_/A vssd1 vssd1 vccd1 vccd1 _3886_/A sky130_fd_sc_hd__o21a_1
X_5623_ _5895_/A vssd1 vssd1 vccd1 vccd1 _5623_/Y sky130_fd_sc_hd__inv_2
X_5554_ _5554_/A _5554_/B vssd1 vssd1 vccd1 vccd1 _5556_/C sky130_fd_sc_hd__xor2_1
X_4505_ _4505_/A _4505_/B vssd1 vssd1 vccd1 vccd1 _4609_/A sky130_fd_sc_hd__nor2_1
X_5485_ _5485_/A _5540_/B vssd1 vssd1 vccd1 vccd1 _5542_/B sky130_fd_sc_hd__and2_1
X_4436_ _4436_/A _4436_/B vssd1 vssd1 vccd1 vccd1 _4548_/B sky130_fd_sc_hd__xnor2_4
X_7224_ _7224_/CLK _7224_/D vssd1 vssd1 vccd1 vccd1 hold75/A sky130_fd_sc_hd__dfxtp_1
X_7155_ _7225_/CLK _7155_/D vssd1 vssd1 vccd1 vccd1 _7155_/Q sky130_fd_sc_hd__dfxtp_1
X_4367_ _4367_/A _3798_/A vssd1 vssd1 vccd1 vccd1 _4367_/X sky130_fd_sc_hd__or2b_1
X_6106_ _6106_/A _6106_/B vssd1 vssd1 vccd1 vccd1 _6108_/A sky130_fd_sc_hd__nand2_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7285__78 vssd1 vssd1 vccd1 vccd1 _7285__78/HI _7393_/A sky130_fd_sc_hd__conb_1
X_7086_ _7099_/A vssd1 vssd1 vccd1 vccd1 _7086_/X sky130_fd_sc_hd__clkbuf_2
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4298_ _5011_/A _5827_/A _4374_/A vssd1 vssd1 vccd1 vccd1 _4298_/Y sky130_fd_sc_hd__o21ai_1
X_6037_ _6037_/A _6133_/B vssd1 vssd1 vccd1 vccd1 _6038_/B sky130_fd_sc_hd__xor2_4
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6939_ _7117_/A vssd1 vssd1 vccd1 vccd1 _6939_/X sky130_fd_sc_hd__clkbuf_2
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5270_ _5271_/A _5271_/B vssd1 vssd1 vccd1 vccd1 _5386_/B sky130_fd_sc_hd__nor2_1
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4221_ _7163_/Q _4572_/A vssd1 vssd1 vccd1 vccd1 _5972_/C sky130_fd_sc_hd__xnor2_4
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4152_ _4553_/A _5017_/A _4152_/C _5016_/A vssd1 vssd1 vccd1 vccd1 _4159_/A sky130_fd_sc_hd__or4b_1
X_4083_ _4083_/A _4083_/B vssd1 vssd1 vccd1 vccd1 _4084_/B sky130_fd_sc_hd__and2_1
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4985_ _7215_/Q vssd1 vssd1 vccd1 vccd1 _5275_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3936_ _7213_/Q _5292_/A vssd1 vssd1 vccd1 vccd1 _3936_/X sky130_fd_sc_hd__and2_1
X_6724_ _6724_/A _6724_/B vssd1 vssd1 vccd1 vccd1 _6730_/B sky130_fd_sc_hd__or2_1
X_3867_ _3867_/A _3867_/B vssd1 vssd1 vccd1 vccd1 _3908_/A sky130_fd_sc_hd__xnor2_1
X_6655_ _6973_/A _6655_/B vssd1 vssd1 vccd1 vccd1 _6656_/B sky130_fd_sc_hd__and2_1
X_5606_ _6539_/A _5606_/B vssd1 vssd1 vccd1 vccd1 _5607_/B sky130_fd_sc_hd__nor2_1
X_6586_ _6586_/A _6586_/B vssd1 vssd1 vccd1 vccd1 _6639_/A sky130_fd_sc_hd__xnor2_2
X_3798_ _3798_/A _4367_/A vssd1 vssd1 vccd1 vccd1 _4339_/A sky130_fd_sc_hd__xnor2_2
XFILLER_11_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5537_ _5515_/A _5537_/B vssd1 vssd1 vccd1 vccd1 _5556_/B sky130_fd_sc_hd__and2b_1
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7207_ _7222_/CLK _7207_/D vssd1 vssd1 vccd1 vccd1 hold83/A sky130_fd_sc_hd__dfxtp_1
X_5468_ _5468_/A _5468_/B vssd1 vssd1 vccd1 vccd1 _5468_/X sky130_fd_sc_hd__or2_1
X_4419_ _4407_/A _4407_/B _4407_/C vssd1 vssd1 vccd1 vccd1 _4495_/A sky130_fd_sc_hd__o21a_1
XFILLER_59_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5399_ _5399_/A _5399_/B vssd1 vssd1 vccd1 vccd1 _5402_/A sky130_fd_sc_hd__xnor2_1
XFILLER_101_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7138_ _7151_/CLK hold18/X vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__dfxtp_1
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7069_ _4400_/A _7062_/X _7068_/X _7060_/X vssd1 vssd1 vccd1 vccd1 _7204_/D sky130_fd_sc_hd__o211a_1
XFILLER_39_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput19 la1_data_in[0] vssd1 vssd1 vccd1 vccd1 _6907_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_52_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4770_ _4770_/A _4770_/B vssd1 vssd1 vccd1 vccd1 _4771_/B sky130_fd_sc_hd__and2_1
XFILLER_60_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3721_ _3721_/A vssd1 vssd1 vccd1 vccd1 _3721_/Y sky130_fd_sc_hd__inv_2
X_6440_ _6432_/B _6432_/C _6022_/A vssd1 vssd1 vccd1 vccd1 _6441_/D sky130_fd_sc_hd__a21oi_1
X_3652_ _3653_/A vssd1 vssd1 vccd1 vccd1 _3652_/Y sky130_fd_sc_hd__inv_2
X_6371_ _6371_/A _6371_/B vssd1 vssd1 vccd1 vccd1 _6374_/A sky130_fd_sc_hd__xnor2_1
X_5322_ _5322_/A _5322_/B vssd1 vssd1 vccd1 vccd1 _5360_/A sky130_fd_sc_hd__nor2_1
XFILLER_88_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5253_ _5253_/A _5253_/B vssd1 vssd1 vccd1 vccd1 _5256_/A sky130_fd_sc_hd__xor2_4
X_4204_ _4216_/A _4204_/B vssd1 vssd1 vccd1 vccd1 _4220_/A sky130_fd_sc_hd__xnor2_1
X_5184_ _4998_/A _4998_/B _5183_/X vssd1 vssd1 vccd1 vccd1 _5361_/B sky130_fd_sc_hd__o21ai_2
XFILLER_56_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4135_ _4279_/A vssd1 vssd1 vccd1 vccd1 _5168_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_95_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7255__48 vssd1 vssd1 vccd1 vccd1 _7255__48/HI _7354_/A sky130_fd_sc_hd__conb_1
X_4066_ _7154_/Q vssd1 vssd1 vccd1 vccd1 _6494_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_56_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4968_ _7215_/Q vssd1 vssd1 vccd1 vccd1 _5133_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4899_ _4899_/A _4899_/B vssd1 vssd1 vccd1 vccd1 _4899_/Y sky130_fd_sc_hd__nor2_1
X_3919_ _4252_/A _3848_/Y _3857_/Y vssd1 vssd1 vccd1 vccd1 _3920_/B sky130_fd_sc_hd__o21ba_1
X_6707_ _6707_/A _6707_/B vssd1 vssd1 vccd1 vccd1 _6707_/X sky130_fd_sc_hd__xor2_2
X_6638_ _6651_/A _6651_/B _6652_/B _6637_/X vssd1 vssd1 vccd1 vccd1 _6640_/A sky130_fd_sc_hd__a31oi_4
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6569_ _6569_/A _6569_/B vssd1 vssd1 vccd1 vccd1 _6592_/B sky130_fd_sc_hd__nand2_1
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5940_ _6947_/A _5953_/A _5953_/B _4328_/B vssd1 vssd1 vccd1 vccd1 _6007_/A sky130_fd_sc_hd__or4b_2
XFILLER_53_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5871_ _5871_/A _5871_/B vssd1 vssd1 vccd1 vccd1 _5879_/A sky130_fd_sc_hd__xnor2_1
X_4822_ _7038_/A _4822_/B _4822_/C vssd1 vssd1 vccd1 vccd1 _4872_/A sky130_fd_sc_hd__nand3_2
XFILLER_33_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4753_ _4748_/A _4790_/A _4790_/B _4752_/Y vssd1 vssd1 vccd1 vccd1 _4757_/B sky130_fd_sc_hd__o31a_1
X_3704_ _3710_/A vssd1 vssd1 vccd1 vccd1 _3709_/A sky130_fd_sc_hd__buf_12
X_4684_ _4684_/A vssd1 vssd1 vccd1 vccd1 _4684_/Y sky130_fd_sc_hd__clkinv_2
X_6423_ _6423_/A _6423_/B vssd1 vssd1 vccd1 vccd1 _6423_/Y sky130_fd_sc_hd__nand2_1
X_3635_ _3635_/A vssd1 vssd1 vccd1 vccd1 _3635_/Y sky130_fd_sc_hd__inv_2
X_6354_ _6354_/A _6309_/A vssd1 vssd1 vccd1 vccd1 _6354_/X sky130_fd_sc_hd__or2b_1
X_6285_ _6285_/A _6342_/A vssd1 vssd1 vccd1 vccd1 _6297_/A sky130_fd_sc_hd__xnor2_2
X_5305_ _5409_/B _5305_/B vssd1 vssd1 vccd1 vccd1 _5307_/B sky130_fd_sc_hd__and2_1
XFILLER_88_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5236_ _5087_/B _5236_/B vssd1 vssd1 vccd1 vccd1 _5236_/X sky130_fd_sc_hd__and2b_1
XFILLER_84_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5167_ _5167_/A vssd1 vssd1 vccd1 vccd1 _5804_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_83_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5098_ _5098_/A _5098_/B vssd1 vssd1 vccd1 vccd1 _5098_/Y sky130_fd_sc_hd__nor2_1
X_4118_ _4382_/B _4118_/B vssd1 vssd1 vccd1 vccd1 _4202_/B sky130_fd_sc_hd__nor2_2
XFILLER_83_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4049_ _6484_/B hold96/A vssd1 vssd1 vccd1 vccd1 _4076_/B sky130_fd_sc_hd__and2b_1
XFILLER_71_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_47_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6070_ _6070_/A _6070_/B _6070_/C vssd1 vssd1 vccd1 vccd1 _6071_/B sky130_fd_sc_hd__nand3_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5021_ _5021_/A _6016_/A vssd1 vssd1 vccd1 vccd1 _5023_/B sky130_fd_sc_hd__xnor2_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6972_ _6693_/A _6964_/X _6971_/X _6967_/X vssd1 vssd1 vccd1 vccd1 _7168_/D sky130_fd_sc_hd__o211a_1
X_5923_ _5923_/A _5923_/B vssd1 vssd1 vccd1 vccd1 _5942_/A sky130_fd_sc_hd__nand2_1
XFILLER_61_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5854_ _5854_/A vssd1 vssd1 vccd1 vccd1 _6560_/A sky130_fd_sc_hd__clkbuf_2
X_4805_ _4819_/A _4805_/B vssd1 vssd1 vccd1 vccd1 _4806_/B sky130_fd_sc_hd__and2_1
X_5785_ _6286_/B _5785_/B vssd1 vssd1 vccd1 vccd1 _5787_/C sky130_fd_sc_hd__nand2_1
X_4736_ _4771_/A _4736_/B vssd1 vssd1 vccd1 vccd1 _4737_/B sky130_fd_sc_hd__or2_1
X_4667_ _4914_/B vssd1 vssd1 vccd1 vccd1 _4674_/A sky130_fd_sc_hd__inv_2
X_7386_ _7386_/A _3677_/Y vssd1 vssd1 vccd1 vccd1 io_out[28] sky130_fd_sc_hd__ebufn_8
X_3618_ _3622_/A vssd1 vssd1 vccd1 vccd1 _3618_/Y sky130_fd_sc_hd__inv_2
X_6406_ _5594_/X hold108/X _6403_/Y _6404_/X _6405_/X vssd1 vssd1 vccd1 vccd1 hold44/A
+ sky130_fd_sc_hd__o221a_1
X_4598_ _4600_/A _4600_/B _4597_/Y vssd1 vssd1 vccd1 vccd1 _4636_/A sky130_fd_sc_hd__o21ai_1
X_6337_ _6280_/A _6280_/B _6336_/X vssd1 vssd1 vccd1 vccd1 _6338_/B sky130_fd_sc_hd__o21a_1
XFILLER_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6268_ _6269_/A _6854_/A vssd1 vssd1 vccd1 vccd1 _6268_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6199_ _6108_/A _6108_/B _6115_/B vssd1 vssd1 vccd1 vccd1 _6199_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_29_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5219_ _5219_/A _5341_/C vssd1 vssd1 vccd1 vccd1 _5222_/A sky130_fd_sc_hd__xnor2_1
XFILLER_17_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5570_ _5570_/A _5570_/B vssd1 vssd1 vccd1 vccd1 _5570_/Y sky130_fd_sc_hd__nor2_1
X_4521_ _4599_/A _4599_/B _4520_/Y vssd1 vssd1 vccd1 vccd1 _4522_/B sky130_fd_sc_hd__a21o_1
X_4452_ _4469_/B _4452_/B vssd1 vssd1 vccd1 vccd1 _4555_/A sky130_fd_sc_hd__xnor2_1
XFILLER_7_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4383_ _4383_/A _4383_/B vssd1 vssd1 vccd1 vccd1 _4384_/B sky130_fd_sc_hd__nor2_1
X_7171_ _7183_/CLK _7171_/D vssd1 vssd1 vccd1 vccd1 _7171_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6122_ _6122_/A _6122_/B vssd1 vssd1 vccd1 vccd1 _6124_/B sky130_fd_sc_hd__xnor2_1
XFILLER_85_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ _6264_/A _6824_/A _5706_/B _5709_/B vssd1 vssd1 vccd1 vccd1 _6054_/B sky130_fd_sc_hd__a31o_1
XFILLER_85_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _5606_/B _5611_/C _4138_/B vssd1 vssd1 vccd1 vccd1 _5004_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6955_ _6480_/A _6949_/X _6954_/X _6952_/X vssd1 vssd1 vccd1 vccd1 _7162_/D sky130_fd_sc_hd__o211a_1
X_5906_ _5932_/A _5931_/A vssd1 vssd1 vccd1 vccd1 _5941_/A sky130_fd_sc_hd__xnor2_1
X_6886_ _6886_/A _6886_/B _6886_/C _6886_/D vssd1 vssd1 vccd1 vccd1 _6887_/C sky130_fd_sc_hd__or4_1
X_5837_ _5870_/A _5870_/B _5836_/X vssd1 vssd1 vccd1 vccd1 _5841_/B sky130_fd_sc_hd__a21o_1
XFILLER_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5768_ _5717_/A _5827_/B _5767_/X vssd1 vssd1 vccd1 vccd1 _5770_/B sky130_fd_sc_hd__a21oi_1
X_4719_ _4948_/A _4948_/B vssd1 vssd1 vccd1 vccd1 _4942_/A sky130_fd_sc_hd__xnor2_1
XFILLER_30_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5699_ _5699_/A _5699_/B vssd1 vssd1 vccd1 vccd1 _5700_/B sky130_fd_sc_hd__xor2_4
XFILLER_30_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7369_ _7369_/A _3657_/Y vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__ebufn_8
XFILLER_1_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6740_ _6740_/A _6740_/B vssd1 vssd1 vccd1 vccd1 _6778_/C sky130_fd_sc_hd__xor2_1
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3952_ hold94/A _4036_/A vssd1 vssd1 vccd1 vccd1 _3960_/A sky130_fd_sc_hd__nand2_1
XFILLER_50_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3883_ _4986_/B _3883_/B vssd1 vssd1 vccd1 vccd1 _3887_/A sky130_fd_sc_hd__or2_1
X_6671_ _6671_/A _6671_/B vssd1 vssd1 vccd1 vccd1 _6672_/B sky130_fd_sc_hd__and2_1
X_5622_ _5756_/A _5897_/B vssd1 vssd1 vccd1 vccd1 _5812_/B sky130_fd_sc_hd__xnor2_4
X_5553_ _5553_/A _5553_/B vssd1 vssd1 vccd1 vccd1 _5554_/B sky130_fd_sc_hd__xnor2_1
X_4504_ _4504_/A _4504_/B vssd1 vssd1 vccd1 vccd1 _4505_/B sky130_fd_sc_hd__and2_1
X_5484_ _6945_/A _5483_/C _6129_/A vssd1 vssd1 vccd1 vccd1 _5540_/B sky130_fd_sc_hd__o21ai_1
X_7223_ _7225_/CLK _7223_/D vssd1 vssd1 vccd1 vccd1 _7223_/Q sky130_fd_sc_hd__dfxtp_1
X_4435_ _4332_/Y _4435_/B vssd1 vssd1 vccd1 vccd1 _4436_/B sky130_fd_sc_hd__and2b_1
X_7154_ _7225_/CLK _7154_/D vssd1 vssd1 vccd1 vccd1 _7154_/Q sky130_fd_sc_hd__dfxtp_1
X_4366_ _4366_/A _4366_/B vssd1 vssd1 vccd1 vccd1 _4949_/A sky130_fd_sc_hd__xnor2_4
XFILLER_98_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6105_ _5262_/X _6102_/X hold126/X _7226_/D vssd1 vssd1 vccd1 vccd1 _7129_/D sky130_fd_sc_hd__o211a_1
XFILLER_98_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7085_ _7085_/A _7093_/B vssd1 vssd1 vccd1 vccd1 _7085_/Y sky130_fd_sc_hd__nand2_1
XFILLER_86_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4297_ _5750_/B _4232_/B _4296_/Y vssd1 vssd1 vccd1 vccd1 _4301_/A sky130_fd_sc_hd__o21ai_2
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _6034_/A _5681_/B _6035_/X vssd1 vssd1 vccd1 vccd1 _6133_/B sky130_fd_sc_hd__a21o_1
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6938_ _6938_/A _6956_/B vssd1 vssd1 vccd1 vccd1 _6938_/Y sky130_fd_sc_hd__nand2_1
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6869_ _6869_/A _6869_/B _6869_/C vssd1 vssd1 vccd1 vccd1 _6869_/X sky130_fd_sc_hd__or3_1
XFILLER_22_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4220_ _4220_/A _4220_/B vssd1 vssd1 vccd1 vccd1 _4421_/A sky130_fd_sc_hd__xnor2_1
XFILLER_95_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4151_ _6439_/A vssd1 vssd1 vccd1 vccd1 _4553_/A sky130_fd_sc_hd__buf_2
XFILLER_95_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4082_ _4083_/A _4083_/B vssd1 vssd1 vccd1 vccd1 _4084_/A sky130_fd_sc_hd__nor2_1
XFILLER_95_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4984_ _6455_/A vssd1 vssd1 vccd1 vccd1 _5287_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_51_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3935_ _4426_/A vssd1 vssd1 vccd1 vccd1 _5292_/A sky130_fd_sc_hd__clkbuf_2
X_6723_ _6723_/A _6723_/B vssd1 vssd1 vccd1 vccd1 _6740_/A sky130_fd_sc_hd__nor2_1
XFILLER_23_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6654_ _6654_/A _6654_/B vssd1 vssd1 vccd1 vccd1 _6667_/A sky130_fd_sc_hd__nand2_1
X_7309__102 vssd1 vssd1 vccd1 vccd1 _7309__102/HI _7417_/A sky130_fd_sc_hd__conb_1
X_3866_ _3910_/A _3998_/B _3865_/X vssd1 vssd1 vccd1 vccd1 _3867_/B sky130_fd_sc_hd__a21oi_1
X_5605_ _6986_/A _5605_/B vssd1 vssd1 vccd1 vccd1 _5802_/A sky130_fd_sc_hd__nor2_1
X_6585_ _6585_/A _6585_/B vssd1 vssd1 vccd1 vccd1 _6611_/A sky130_fd_sc_hd__xor2_1
X_3797_ _4285_/A _3797_/B vssd1 vssd1 vccd1 vccd1 _4367_/A sky130_fd_sc_hd__xnor2_2
X_5536_ _5529_/A _5529_/B _5530_/A vssd1 vssd1 vccd1 vccd1 _5569_/A sky130_fd_sc_hd__a21o_1
X_5467_ _5528_/A _5467_/B vssd1 vssd1 vccd1 vccd1 _5475_/A sky130_fd_sc_hd__xnor2_1
X_4418_ _4418_/A vssd1 vssd1 vccd1 vccd1 _4496_/B sky130_fd_sc_hd__inv_2
X_7206_ _7222_/CLK _7206_/D vssd1 vssd1 vccd1 vccd1 hold85/A sky130_fd_sc_hd__dfxtp_1
X_5398_ _5398_/A _5490_/B vssd1 vssd1 vccd1 vccd1 _5399_/B sky130_fd_sc_hd__nor2_1
X_7137_ _7224_/CLK hold42/X vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__dfxtp_1
X_4349_ _5604_/A _7171_/Q vssd1 vssd1 vccd1 vccd1 _5190_/A sky130_fd_sc_hd__nor2_1
X_7068_ hold87/X _7091_/B vssd1 vssd1 vccd1 vccd1 _7068_/X sky130_fd_sc_hd__or2_1
X_6019_ _6266_/B _6019_/B vssd1 vssd1 vccd1 vccd1 _6106_/A sky130_fd_sc_hd__nand2_1
XFILLER_100_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3720_ _3721_/A vssd1 vssd1 vccd1 vccd1 _3720_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3651_ _3653_/A vssd1 vssd1 vccd1 vccd1 _3651_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6370_ _6990_/A _6370_/B vssd1 vssd1 vccd1 vccd1 _6371_/B sky130_fd_sc_hd__xnor2_1
X_5321_ _5321_/A _5321_/B _5321_/C vssd1 vssd1 vccd1 vccd1 _5322_/B sky130_fd_sc_hd__nor3_1
XFILLER_88_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5252_ _5372_/A _5372_/B vssd1 vssd1 vccd1 vccd1 _5253_/B sky130_fd_sc_hd__xnor2_4
X_4203_ _4342_/A _4342_/B vssd1 vssd1 vccd1 vccd1 _4236_/A sky130_fd_sc_hd__xnor2_4
X_5183_ _5183_/A _5183_/B vssd1 vssd1 vccd1 vccd1 _5183_/X sky130_fd_sc_hd__or2_1
XFILLER_3_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4134_ _4375_/B _4134_/B vssd1 vssd1 vccd1 vccd1 _4149_/A sky130_fd_sc_hd__xor2_1
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4065_ _4065_/A _4065_/B vssd1 vssd1 vccd1 vccd1 _4083_/A sky130_fd_sc_hd__xnor2_1
XFILLER_36_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4967_ _5145_/A _5145_/B vssd1 vssd1 vccd1 vccd1 _4972_/A sky130_fd_sc_hd__nor2_1
XFILLER_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4898_ _4902_/A _4898_/B vssd1 vssd1 vccd1 vccd1 _4919_/B sky130_fd_sc_hd__and2b_1
X_3918_ _3918_/A _3966_/A vssd1 vssd1 vccd1 vccd1 _4019_/A sky130_fd_sc_hd__xnor2_2
X_6706_ _6706_/A _6706_/B _6706_/C _6705_/X vssd1 vssd1 vccd1 vccd1 _6707_/B sky130_fd_sc_hd__or4b_4
X_3849_ _7185_/Q vssd1 vssd1 vccd1 vccd1 _4526_/B sky130_fd_sc_hd__clkbuf_2
X_6637_ _6636_/B _6637_/B vssd1 vssd1 vccd1 vccd1 _6637_/X sky130_fd_sc_hd__and2b_1
X_6568_ _6981_/A _6568_/B vssd1 vssd1 vccd1 vccd1 _6569_/B sky130_fd_sc_hd__nand2_1
XFILLER_3_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5519_ _5456_/A _5456_/B _5518_/X vssd1 vssd1 vccd1 vccd1 _5520_/B sky130_fd_sc_hd__a21boi_1
X_6499_ _6506_/A vssd1 vssd1 vccd1 vccd1 _6520_/B sky130_fd_sc_hd__clkinv_2
XFILLER_3_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5870_ _5870_/A _5870_/B vssd1 vssd1 vccd1 vccd1 _5883_/A sky130_fd_sc_hd__xnor2_2
XFILLER_18_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4821_ _4821_/A _4821_/B vssd1 vssd1 vccd1 vccd1 _4822_/C sky130_fd_sc_hd__or2_1
XFILLER_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4752_ _4808_/A _4808_/B vssd1 vssd1 vccd1 vccd1 _4752_/Y sky130_fd_sc_hd__nand2_1
X_4683_ _4838_/A _4593_/B _4838_/B _4682_/Y vssd1 vssd1 vccd1 vccd1 _4739_/B sky130_fd_sc_hd__o31a_1
X_3703_ _3703_/A vssd1 vssd1 vccd1 vccd1 _3703_/Y sky130_fd_sc_hd__inv_2
X_3634_ _3635_/A vssd1 vssd1 vccd1 vccd1 _3634_/Y sky130_fd_sc_hd__inv_2
X_6422_ _6423_/A _6423_/B vssd1 vssd1 vccd1 vccd1 _6424_/A sky130_fd_sc_hd__nor2_1
X_6353_ _6353_/A _6353_/B vssd1 vssd1 vccd1 vccd1 _6356_/A sky130_fd_sc_hd__xor2_1
XFILLER_88_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6284_ _6219_/A _6219_/B _6283_/X vssd1 vssd1 vccd1 vccd1 _6342_/A sky130_fd_sc_hd__o21a_1
X_5304_ _5606_/B _5304_/B vssd1 vssd1 vccd1 vccd1 _5305_/B sky130_fd_sc_hd__or2_1
XFILLER_88_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5235_ _5354_/B _5235_/B vssd1 vssd1 vccd1 vccd1 _5238_/A sky130_fd_sc_hd__xnor2_1
XFILLER_96_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5166_ _6850_/A _5166_/B vssd1 vssd1 vccd1 vccd1 _5178_/A sky130_fd_sc_hd__xor2_2
XFILLER_56_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5097_ _5098_/A _5098_/B vssd1 vssd1 vccd1 vccd1 _5097_/Y sky130_fd_sc_hd__nand2_1
X_4117_ _4117_/A _4117_/B vssd1 vssd1 vccd1 vccd1 _4118_/B sky130_fd_sc_hd__and2_1
XFILLER_83_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4048_ _7155_/Q vssd1 vssd1 vccd1 vccd1 _6484_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_56_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5999_ _5980_/B _5999_/B vssd1 vssd1 vccd1 vccd1 _6000_/A sky130_fd_sc_hd__and2b_1
XFILLER_33_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5020_ _6449_/A vssd1 vssd1 vccd1 vccd1 _6464_/A sky130_fd_sc_hd__clkbuf_2
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6971_ _6971_/A _6975_/B vssd1 vssd1 vccd1 vccd1 _6971_/X sky130_fd_sc_hd__or2_1
XFILLER_80_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5922_ _5922_/A _5938_/A vssd1 vssd1 vccd1 vccd1 _5923_/B sky130_fd_sc_hd__or2_1
X_5853_ _6301_/A _6174_/A _6241_/A _6061_/B vssd1 vssd1 vccd1 vccd1 _5856_/A sky130_fd_sc_hd__o211a_1
X_4804_ _4819_/A _4805_/B vssd1 vssd1 vccd1 vccd1 _4806_/A sky130_fd_sc_hd__nor2_1
X_5784_ _5784_/A _5784_/B vssd1 vssd1 vccd1 vccd1 _5785_/B sky130_fd_sc_hd__nand2_1
XFILLER_34_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4735_ _4771_/A _4736_/B vssd1 vssd1 vccd1 vccd1 _4737_/A sky130_fd_sc_hd__nand2_1
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4666_ _4666_/A _4666_/B vssd1 vssd1 vccd1 vccd1 _4723_/A sky130_fd_sc_hd__nor2_1
X_4597_ _4597_/A _4597_/B vssd1 vssd1 vccd1 vccd1 _4597_/Y sky130_fd_sc_hd__nand2_1
X_3617_ _3742_/A vssd1 vssd1 vccd1 vccd1 _3622_/A sky130_fd_sc_hd__buf_12
X_7385_ _7385_/A _3676_/Y vssd1 vssd1 vccd1 vccd1 io_out[27] sky130_fd_sc_hd__ebufn_8
X_6405_ _7099_/A vssd1 vssd1 vccd1 vccd1 _6405_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_1_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6336_ _6336_/A _6282_/B vssd1 vssd1 vccd1 vccd1 _6336_/X sky130_fd_sc_hd__or2b_1
XFILLER_88_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6267_ _6199_/Y _6266_/Y _5143_/X vssd1 vssd1 vccd1 vccd1 _6854_/A sky130_fd_sc_hd__a21o_2
XFILLER_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6198_ _6198_/A _6198_/B vssd1 vssd1 vccd1 vccd1 _6213_/A sky130_fd_sc_hd__or2_1
X_5218_ _5218_/A _5218_/B vssd1 vssd1 vccd1 vccd1 _5341_/C sky130_fd_sc_hd__xor2_1
XFILLER_69_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5149_ _5149_/A _5149_/B vssd1 vssd1 vccd1 vccd1 _5150_/B sky130_fd_sc_hd__nor2_1
XFILLER_84_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4520_ _4520_/A _4520_/B vssd1 vssd1 vccd1 vccd1 _4520_/Y sky130_fd_sc_hd__nor2_1
X_4451_ _5644_/A _4567_/B vssd1 vssd1 vccd1 vccd1 _4666_/A sky130_fd_sc_hd__and2_1
XFILLER_7_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7170_ _7172_/CLK _7170_/D vssd1 vssd1 vccd1 vccd1 _7170_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4382_ _4382_/A _4382_/B _4382_/C vssd1 vssd1 vccd1 vccd1 _4383_/B sky130_fd_sc_hd__nor3_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6121_ _6121_/A _6206_/B vssd1 vssd1 vccd1 vccd1 _6122_/B sky130_fd_sc_hd__or2_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6052_ _6531_/A vssd1 vssd1 vccd1 vccd1 _6824_/A sky130_fd_sc_hd__clkbuf_2
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _5168_/A vssd1 vssd1 vccd1 vccd1 _5611_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_66_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6954_ _6954_/A _6954_/B vssd1 vssd1 vccd1 vccd1 _6954_/X sky130_fd_sc_hd__or2_1
X_5905_ _5914_/A _5914_/B _5902_/B _5923_/A vssd1 vssd1 vccd1 vccd1 _5931_/A sky130_fd_sc_hd__o31a_1
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6885_ hold23/X _3750_/X _5595_/X _6884_/Y vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__o211a_1
X_5836_ _5835_/B _5836_/B vssd1 vssd1 vccd1 vccd1 _5836_/X sky130_fd_sc_hd__and2b_1
X_5767_ _7019_/A _6480_/A vssd1 vssd1 vccd1 vccd1 _5767_/X sky130_fd_sc_hd__and2_1
X_4718_ _4936_/A _4936_/B _4717_/Y vssd1 vssd1 vccd1 vccd1 _4948_/B sky130_fd_sc_hd__a21oi_1
X_5698_ _5698_/A _5698_/B vssd1 vssd1 vccd1 vccd1 _5700_/A sky130_fd_sc_hd__nand2_2
X_4649_ _4649_/A _4649_/B vssd1 vssd1 vccd1 vccd1 _4702_/C sky130_fd_sc_hd__nor2_1
X_7368_ _7368_/A _3656_/Y vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__ebufn_8
X_6319_ _6319_/A _6319_/B vssd1 vssd1 vccd1 vccd1 _6319_/X sky130_fd_sc_hd__xor2_2
XFILLER_39_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3951_ _4208_/A _7215_/Q vssd1 vssd1 vccd1 vccd1 _4036_/A sky130_fd_sc_hd__or2b_1
XFILLER_16_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6670_ _6671_/A _6671_/B vssd1 vssd1 vccd1 vccd1 _6672_/A sky130_fd_sc_hd__nor2_1
X_3882_ _5274_/A _4411_/A vssd1 vssd1 vccd1 vccd1 _3883_/B sky130_fd_sc_hd__nor2_1
XFILLER_31_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5621_ _5787_/A _5737_/C _5985_/B vssd1 vssd1 vccd1 vccd1 _5897_/B sky130_fd_sc_hd__a21o_2
X_5552_ _5552_/A _5552_/B vssd1 vssd1 vccd1 vccd1 _5553_/B sky130_fd_sc_hd__nor2_1
X_4503_ _4506_/A _4506_/B vssd1 vssd1 vccd1 vccd1 _4503_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5483_ _6129_/A _6945_/A _5483_/C vssd1 vssd1 vccd1 vccd1 _5485_/A sky130_fd_sc_hd__or3_1
X_4434_ _4437_/A _4437_/B vssd1 vssd1 vccd1 vccd1 _4548_/A sky130_fd_sc_hd__xnor2_2
X_7222_ _7222_/CLK _7222_/D vssd1 vssd1 vccd1 vccd1 hold96/A sky130_fd_sc_hd__dfxtp_1
X_7153_ _7225_/CLK _7153_/D vssd1 vssd1 vccd1 vccd1 _7153_/Q sky130_fd_sc_hd__dfxtp_2
X_4365_ _5218_/A _5073_/B vssd1 vssd1 vccd1 vccd1 _4366_/B sky130_fd_sc_hd__xor2_4
X_7084_ hold91/X _7075_/X _7083_/Y _7073_/X vssd1 vssd1 vccd1 vccd1 hold92/A sky130_fd_sc_hd__o211a_1
X_6104_ _6391_/A hold32/X vssd1 vssd1 vccd1 vccd1 _6104_/X sky130_fd_sc_hd__or2_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6035_ _6035_/A _6035_/B vssd1 vssd1 vccd1 vccd1 _6035_/X sky130_fd_sc_hd__and2_1
X_4296_ _6713_/A _4296_/B vssd1 vssd1 vccd1 vccd1 _4296_/Y sky130_fd_sc_hd__nand2_1
XFILLER_100_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6937_ _7080_/A vssd1 vssd1 vccd1 vccd1 _6956_/B sky130_fd_sc_hd__clkbuf_2
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6868_ _6869_/A _6869_/B _6869_/C vssd1 vssd1 vccd1 vccd1 _6877_/B sky130_fd_sc_hd__o21ai_1
XFILLER_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5819_ _5818_/B _5819_/B vssd1 vssd1 vccd1 vccd1 _5820_/B sky130_fd_sc_hd__and2b_1
X_6799_ _6799_/A _6799_/B vssd1 vssd1 vccd1 vccd1 _6824_/B sky130_fd_sc_hd__and2_1
XFILLER_10_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7276__69 vssd1 vssd1 vccd1 vccd1 _7276__69/HI _7375_/A sky130_fd_sc_hd__conb_1
XFILLER_92_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4150_ _4150_/A _4150_/B vssd1 vssd1 vccd1 vccd1 _4164_/A sky130_fd_sc_hd__nand2_2
XFILLER_95_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4081_ _4216_/A _4204_/B _4080_/Y vssd1 vssd1 vccd1 vccd1 _4083_/B sky130_fd_sc_hd__o21a_1
XFILLER_95_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7290__83 vssd1 vssd1 vccd1 vccd1 _7290__83/HI _7398_/A sky130_fd_sc_hd__conb_1
XFILLER_36_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4983_ _6470_/A vssd1 vssd1 vccd1 vccd1 _6455_/A sky130_fd_sc_hd__buf_2
X_3934_ _7213_/Q _7212_/Q vssd1 vssd1 vccd1 vccd1 _3944_/B sky130_fd_sc_hd__xor2_4
X_6722_ _6722_/A _6722_/B vssd1 vssd1 vccd1 vccd1 _6723_/B sky130_fd_sc_hd__nor2_1
X_6653_ _6947_/A _6653_/B vssd1 vssd1 vccd1 vccd1 _6654_/B sky130_fd_sc_hd__nand2_1
X_3865_ _7196_/Q _4392_/B vssd1 vssd1 vccd1 vccd1 _3865_/X sky130_fd_sc_hd__and2_1
X_5604_ _5604_/A vssd1 vssd1 vccd1 vccd1 _6986_/A sky130_fd_sc_hd__clkbuf_2
X_6584_ _6584_/A _6584_/B vssd1 vssd1 vccd1 vccd1 _6585_/B sky130_fd_sc_hd__xnor2_1
X_3796_ _4344_/A _4344_/B vssd1 vssd1 vccd1 vccd1 _3797_/B sky130_fd_sc_hd__xor2_2
X_5535_ _5262_/X _5533_/X hold55/X _7226_/D vssd1 vssd1 vccd1 vccd1 hold57/A sky130_fd_sc_hd__o211a_1
X_5466_ _5466_/A _5527_/A vssd1 vssd1 vccd1 vccd1 _5467_/B sky130_fd_sc_hd__xnor2_1
X_4417_ _4538_/A _4538_/B _4416_/Y _7085_/A vssd1 vssd1 vccd1 vccd1 _4418_/A sky130_fd_sc_hd__o22a_1
X_7205_ _7222_/CLK _7205_/D vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__dfxtp_2
X_5397_ _7096_/A _5397_/B _5397_/C vssd1 vssd1 vccd1 vccd1 _5490_/B sky130_fd_sc_hd__and3_1
XFILLER_98_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7136_ _7224_/CLK hold52/X vssd1 vssd1 vccd1 vccd1 hold51/A sky130_fd_sc_hd__dfxtp_1
X_4348_ _7174_/Q vssd1 vssd1 vccd1 vccd1 _5604_/A sky130_fd_sc_hd__inv_2
XFILLER_100_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7067_ _7043_/A _7062_/X _7066_/Y _7060_/X vssd1 vssd1 vccd1 vccd1 _7203_/D sky130_fd_sc_hd__o211a_1
XFILLER_59_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4279_ _4279_/A _5021_/A vssd1 vssd1 vccd1 vccd1 _4279_/Y sky130_fd_sc_hd__nand2_1
XFILLER_67_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6018_ _7159_/Q _6483_/A vssd1 vssd1 vccd1 vccd1 _6019_/B sky130_fd_sc_hd__or2_1
XFILLER_100_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3650_ _3653_/A vssd1 vssd1 vccd1 vccd1 _3650_/Y sky130_fd_sc_hd__inv_2
X_5320_ _5321_/A _5321_/B _5321_/C vssd1 vssd1 vccd1 vccd1 _5322_/A sky130_fd_sc_hd__o21a_1
X_5251_ _5100_/A _5100_/B _5250_/X vssd1 vssd1 vccd1 vccd1 _5372_/B sky130_fd_sc_hd__o21ai_4
X_4202_ _4202_/A _4202_/B vssd1 vssd1 vccd1 vccd1 _4342_/B sky130_fd_sc_hd__xor2_4
X_5182_ _5265_/A _5265_/B vssd1 vssd1 vccd1 vccd1 _5361_/A sky130_fd_sc_hd__xor2_2
X_4133_ _4133_/A _4133_/B vssd1 vssd1 vccd1 vccd1 _4134_/B sky130_fd_sc_hd__nand2_1
X_4064_ _4064_/A _4064_/B vssd1 vssd1 vccd1 vccd1 _4065_/B sky130_fd_sc_hd__xnor2_1
XFILLER_28_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4966_ _3887_/A _3886_/B _3886_/A vssd1 vssd1 vccd1 vccd1 _4974_/A sky130_fd_sc_hd__o21bai_1
X_6705_ _6673_/X _6703_/X _6672_/A _6704_/X vssd1 vssd1 vccd1 vccd1 _6705_/X sky130_fd_sc_hd__a211o_1
X_4897_ _4882_/A _4847_/B _4910_/A vssd1 vssd1 vccd1 vccd1 _4898_/B sky130_fd_sc_hd__a21bo_1
X_3917_ _3996_/A _3995_/A _3995_/B _3912_/B _3912_/A vssd1 vssd1 vccd1 vccd1 _3966_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_20_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3848_ _4011_/A _3922_/B _5267_/A vssd1 vssd1 vccd1 vccd1 _3848_/Y sky130_fd_sc_hd__a21oi_2
X_6636_ _6637_/B _6636_/B vssd1 vssd1 vccd1 vccd1 _6652_/B sky130_fd_sc_hd__xnor2_2
X_3779_ _7169_/Q vssd1 vssd1 vccd1 vccd1 _5619_/B sky130_fd_sc_hd__clkbuf_2
X_6567_ _6981_/A _6568_/B vssd1 vssd1 vccd1 vccd1 _6569_/A sky130_fd_sc_hd__or2_1
X_5518_ _5518_/A _5457_/A vssd1 vssd1 vccd1 vccd1 _5518_/X sky130_fd_sc_hd__or2b_1
X_6498_ _6493_/X _6505_/A _6487_/X _6497_/Y vssd1 vssd1 vccd1 vccd1 _6506_/A sky130_fd_sc_hd__a211o_1
XFILLER_79_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5449_ _6524_/A vssd1 vssd1 vccd1 vccd1 _6162_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_87_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7119_ _7222_/CLK _7119_/D vssd1 vssd1 vccd1 vccd1 hold93/A sky130_fd_sc_hd__dfxtp_1
XFILLER_59_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7246__39 vssd1 vssd1 vccd1 vccd1 _7246__39/HI _7345_/A sky130_fd_sc_hd__conb_1
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7260__53 vssd1 vssd1 vccd1 vccd1 _7260__53/HI _7359_/A sky130_fd_sc_hd__conb_1
X_4820_ _4820_/A _4820_/B vssd1 vssd1 vccd1 vccd1 _4824_/A sky130_fd_sc_hd__xnor2_2
XFILLER_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4751_ _4838_/B _4751_/B vssd1 vssd1 vccd1 vccd1 _4808_/B sky130_fd_sc_hd__nor2_1
X_4682_ _4593_/B _4838_/B _4838_/A vssd1 vssd1 vccd1 vccd1 _4682_/Y sky130_fd_sc_hd__o21ai_1
X_3702_ _3703_/A vssd1 vssd1 vccd1 vccd1 _3702_/Y sky130_fd_sc_hd__inv_2
X_3633_ _3635_/A vssd1 vssd1 vccd1 vccd1 _3633_/Y sky130_fd_sc_hd__inv_2
X_6421_ _6421_/A _6538_/A vssd1 vssd1 vccd1 vccd1 _6423_/B sky130_fd_sc_hd__xnor2_1
X_6352_ _6385_/B _6352_/B vssd1 vssd1 vccd1 vccd1 _6353_/B sky130_fd_sc_hd__xnor2_1
X_5303_ _6240_/A _5304_/B vssd1 vssd1 vccd1 vccd1 _5409_/B sky130_fd_sc_hd__nand2_1
X_6283_ _6283_/A _6222_/B vssd1 vssd1 vccd1 vccd1 _6283_/X sky130_fd_sc_hd__or2b_1
X_5234_ _5234_/A _5353_/B vssd1 vssd1 vccd1 vccd1 _5235_/B sky130_fd_sc_hd__xor2_1
X_5165_ _5348_/S _5165_/B vssd1 vssd1 vccd1 vccd1 _5166_/B sky130_fd_sc_hd__or2_1
XFILLER_96_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4116_ _4117_/A _4117_/B vssd1 vssd1 vccd1 vccd1 _4382_/B sky130_fd_sc_hd__nor2_1
XFILLER_29_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5096_ _5096_/A _5096_/B vssd1 vssd1 vccd1 vccd1 _5100_/A sky130_fd_sc_hd__xnor2_2
X_4047_ _6016_/A vssd1 vssd1 vccd1 vccd1 _6109_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5998_ _6000_/B _5998_/B _5998_/C vssd1 vssd1 vccd1 vccd1 _5998_/Y sky130_fd_sc_hd__nor3_1
X_4949_ _4949_/A _4369_/B vssd1 vssd1 vccd1 vccd1 _5107_/A sky130_fd_sc_hd__or2b_1
X_6619_ _6619_/A _6619_/B vssd1 vssd1 vccd1 vccd1 _6651_/B sky130_fd_sc_hd__nand2_1
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6970_ _5143_/X _6964_/X _6969_/X _6967_/X vssd1 vssd1 vccd1 vccd1 _7167_/D sky130_fd_sc_hd__o211a_1
XFILLER_53_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5921_ _5924_/A _5924_/B vssd1 vssd1 vccd1 vccd1 _5926_/A sky130_fd_sc_hd__and2b_1
XFILLER_65_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5852_ _6160_/A vssd1 vssd1 vccd1 vccd1 _6241_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4803_ _6933_/A _4803_/B vssd1 vssd1 vccd1 vccd1 _4805_/B sky130_fd_sc_hd__xnor2_1
X_5783_ _5784_/A _5783_/B vssd1 vssd1 vccd1 vccd1 _6286_/B sky130_fd_sc_hd__or2_1
X_4734_ _4734_/A _4734_/B vssd1 vssd1 vccd1 vccd1 _4736_/B sky130_fd_sc_hd__nor2_1
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4665_ _4665_/A _4665_/B vssd1 vssd1 vccd1 vccd1 _4684_/A sky130_fd_sc_hd__xnor2_2
X_4596_ _4586_/A _4586_/B _4587_/B _4663_/A _4663_/B vssd1 vssd1 vccd1 vccd1 _4600_/B
+ sky130_fd_sc_hd__o32a_2
X_7384_ _7384_/A _3675_/Y vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__ebufn_8
X_6404_ _6403_/A _6403_/B _6879_/A vssd1 vssd1 vccd1 vccd1 _6404_/X sky130_fd_sc_hd__a21o_1
X_3616_ _3616_/A vssd1 vssd1 vccd1 vccd1 _3616_/Y sky130_fd_sc_hd__inv_2
X_6335_ _6335_/A _6362_/B vssd1 vssd1 vccd1 vccd1 _6372_/B sky130_fd_sc_hd__xnor2_1
X_6266_ _6943_/A _6266_/B vssd1 vssd1 vccd1 vccd1 _6266_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6197_ _5262_/X _6194_/X _6195_/X _6196_/X vssd1 vssd1 vccd1 vccd1 _7130_/D sky130_fd_sc_hd__o211a_1
X_5217_ _5446_/A _5446_/B vssd1 vssd1 vccd1 vccd1 _5218_/B sky130_fd_sc_hd__xnor2_1
X_5148_ _5148_/A _5148_/B _5148_/C vssd1 vssd1 vccd1 vccd1 _5149_/B sky130_fd_sc_hd__and3_1
XFILLER_56_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5079_ _5690_/A vssd1 vssd1 vccd1 vccd1 _5689_/A sky130_fd_sc_hd__buf_2
XFILLER_44_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7230__23 vssd1 vssd1 vccd1 vccd1 _7230__23/HI _7329_/A sky130_fd_sc_hd__conb_1
XFILLER_31_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4450_ _5026_/A _4450_/B vssd1 vssd1 vccd1 vccd1 _4567_/B sky130_fd_sc_hd__xnor2_2
XFILLER_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4381_ _4382_/A _4382_/B _4382_/C vssd1 vssd1 vccd1 vccd1 _4383_/A sky130_fd_sc_hd__o21a_1
X_6120_ _6120_/A _6120_/B _7025_/A vssd1 vssd1 vccd1 vccd1 _6206_/B sky130_fd_sc_hd__and3_1
XFILLER_98_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6051_ _6154_/A _6154_/B vssd1 vssd1 vccd1 vccd1 _6055_/A sky130_fd_sc_hd__xor2_2
XFILLER_100_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5002_ _5002_/A vssd1 vssd1 vccd1 vccd1 _5606_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6953_ hold123/X _6949_/X _6950_/X _6952_/X vssd1 vssd1 vccd1 vccd1 _7161_/D sky130_fd_sc_hd__o211a_1
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5904_ _5922_/A _5938_/A vssd1 vssd1 vccd1 vccd1 _5923_/A sky130_fd_sc_hd__nand2_1
X_6884_ _6878_/Y _6883_/Y _5113_/X vssd1 vssd1 vccd1 vccd1 _6884_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_41_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5835_ _5836_/B _5835_/B vssd1 vssd1 vccd1 vccd1 _5870_/B sky130_fd_sc_hd__xnor2_1
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5766_ _6466_/B vssd1 vssd1 vccd1 vccd1 _6480_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4717_ _4717_/A _4717_/B vssd1 vssd1 vccd1 vccd1 _4717_/Y sky130_fd_sc_hd__nor2_1
X_5697_ _6140_/A _5719_/B vssd1 vssd1 vccd1 vccd1 _5698_/B sky130_fd_sc_hd__nand2_1
X_4648_ _4730_/A _4730_/B vssd1 vssd1 vccd1 vccd1 _4731_/A sky130_fd_sc_hd__and2_1
XFILLER_89_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4579_ _4579_/A _4579_/B vssd1 vssd1 vccd1 vccd1 _4580_/B sky130_fd_sc_hd__or2_1
X_7367_ _7367_/A _3653_/Y vssd1 vssd1 vccd1 vccd1 io_out[9] sky130_fd_sc_hd__ebufn_8
XFILLER_89_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6318_ _6258_/A _6258_/B _6317_/X vssd1 vssd1 vccd1 vccd1 _6319_/B sky130_fd_sc_hd__a21o_1
X_6249_ _6314_/A _6314_/B vssd1 vssd1 vccd1 vccd1 _6250_/B sky130_fd_sc_hd__xor2_1
XFILLER_84_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3950_ _7220_/Q vssd1 vssd1 vccd1 vccd1 _4208_/A sky130_fd_sc_hd__clkbuf_2
X_3881_ _7211_/Q vssd1 vssd1 vccd1 vccd1 _4411_/A sky130_fd_sc_hd__inv_2
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5620_ _5625_/B vssd1 vssd1 vccd1 vccd1 _5985_/B sky130_fd_sc_hd__clkbuf_2
X_5551_ _5551_/A _5551_/B _5551_/C vssd1 vssd1 vccd1 vccd1 _5552_/B sky130_fd_sc_hd__and3_1
X_4502_ _4502_/A _4763_/A vssd1 vssd1 vccd1 vccd1 _4507_/A sky130_fd_sc_hd__xnor2_1
X_7221_ _7221_/CLK hold95/X vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__dfxtp_1
X_5482_ _6209_/A vssd1 vssd1 vccd1 vccd1 _6264_/A sky130_fd_sc_hd__clkbuf_2
X_4433_ _6475_/A _4550_/A _4659_/A _4641_/A _4429_/A vssd1 vssd1 vccd1 vccd1 _4437_/B
+ sky130_fd_sc_hd__a32oi_4
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7152_ _7225_/CLK _7152_/D vssd1 vssd1 vccd1 vccd1 _7152_/Q sky130_fd_sc_hd__dfxtp_1
X_4364_ _5047_/A _5047_/B vssd1 vssd1 vccd1 vccd1 _5073_/B sky130_fd_sc_hd__xnor2_2
X_7083_ _7083_/A _7093_/B vssd1 vssd1 vccd1 vccd1 _7083_/Y sky130_fd_sc_hd__nand2_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6103_ _6845_/A vssd1 vssd1 vccd1 vccd1 _6391_/A sky130_fd_sc_hd__clkbuf_1
X_4295_ _4374_/A _4375_/B _4289_/A _4289_/B vssd1 vssd1 vccd1 vccd1 _4370_/A sky130_fd_sc_hd__a22o_1
XFILLER_100_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6034_ _6034_/A _6129_/B vssd1 vssd1 vccd1 vccd1 _6037_/A sky130_fd_sc_hd__xnor2_4
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6936_ _7052_/A vssd1 vssd1 vccd1 vccd1 _7080_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6867_ _6873_/A _6873_/B vssd1 vssd1 vccd1 vccd1 _6869_/C sky130_fd_sc_hd__xor2_1
X_6798_ _6797_/A _6797_/B _6797_/C vssd1 vssd1 vccd1 vccd1 _6799_/B sky130_fd_sc_hd__o21ai_1
XFILLER_22_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5818_ _5819_/B _5818_/B vssd1 vssd1 vccd1 vccd1 _5859_/B sky130_fd_sc_hd__and2b_1
X_5749_ _5749_/A vssd1 vssd1 vccd1 vccd1 _6994_/A sky130_fd_sc_hd__buf_2
XFILLER_41_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7419_ _7419_/A _3709_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[23] sky130_fd_sc_hd__ebufn_8
XFILLER_1_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4080_ _4197_/A _4080_/B vssd1 vssd1 vccd1 vccd1 _4080_/Y sky130_fd_sc_hd__nand2_1
XFILLER_76_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4982_ _6109_/A vssd1 vssd1 vccd1 vccd1 _6470_/A sky130_fd_sc_hd__buf_2
X_3933_ _3933_/A _4996_/B vssd1 vssd1 vccd1 vccd1 _3983_/A sky130_fd_sc_hd__xnor2_1
XFILLER_16_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6721_ _6722_/A _6722_/B vssd1 vssd1 vccd1 vccd1 _6723_/A sky130_fd_sc_hd__and2_1
X_3864_ _7195_/Q vssd1 vssd1 vccd1 vccd1 _4392_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6652_ _6652_/A _6652_/B vssd1 vssd1 vccd1 vccd1 _6671_/A sky130_fd_sc_hd__xor2_1
X_5603_ _5643_/B _5603_/B vssd1 vssd1 vccd1 vccd1 _5614_/A sky130_fd_sc_hd__nand2_1
X_3795_ _4355_/A _4354_/A vssd1 vssd1 vccd1 vccd1 _4344_/B sky130_fd_sc_hd__xor2_2
X_6583_ _6583_/A _6745_/A vssd1 vssd1 vccd1 vccd1 _6585_/A sky130_fd_sc_hd__xor2_1
X_5534_ _5594_/A hold56/X vssd1 vssd1 vccd1 vccd1 hold55/A sky130_fd_sc_hd__or2_1
X_5465_ _5367_/A _5367_/B _5464_/X vssd1 vssd1 vccd1 vccd1 _5527_/A sky130_fd_sc_hd__o21a_1
X_4416_ _4540_/B _4416_/B vssd1 vssd1 vccd1 vccd1 _4416_/Y sky130_fd_sc_hd__nand2_1
X_7204_ _7222_/CLK _7204_/D vssd1 vssd1 vccd1 vccd1 _7204_/Q sky130_fd_sc_hd__dfxtp_1
X_7135_ _7151_/CLK hold44/X vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__dfxtp_1
X_5396_ _7096_/A _5397_/B _5397_/C vssd1 vssd1 vccd1 vccd1 _5398_/A sky130_fd_sc_hd__a21oi_1
XFILLER_101_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4347_ _7174_/Q _6563_/A vssd1 vssd1 vccd1 vccd1 _4350_/A sky130_fd_sc_hd__nor2_1
XFILLER_98_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4278_ _5750_/B _4278_/B vssd1 vssd1 vccd1 vccd1 _5826_/A sky130_fd_sc_hd__nand2_4
X_7066_ _7066_/A _7072_/B vssd1 vssd1 vccd1 vccd1 _7066_/Y sky130_fd_sc_hd__nand2_1
X_6017_ _7156_/Q vssd1 vssd1 vccd1 vccd1 _6483_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_74_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6919_ _7116_/A hold46/X vssd1 vssd1 vccd1 vccd1 hold45/A sky130_fd_sc_hd__nor2_1
XFILLER_52_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5250_ _5250_/A _5250_/B vssd1 vssd1 vccd1 vccd1 _5250_/X sky130_fd_sc_hd__or2_1
X_4201_ _4188_/A _4188_/B _4239_/A vssd1 vssd1 vccd1 vccd1 _4342_/A sky130_fd_sc_hd__o21ai_4
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5181_ _5181_/A _5181_/B vssd1 vssd1 vccd1 vccd1 _5265_/B sky130_fd_sc_hd__xor2_1
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4132_ _5784_/B _5688_/A vssd1 vssd1 vccd1 vccd1 _4133_/B sky130_fd_sc_hd__nand2_1
XFILLER_83_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4063_ _5016_/A _6938_/A _4038_/A vssd1 vssd1 vccd1 vccd1 _4064_/B sky130_fd_sc_hd__a21oi_1
XFILLER_83_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4965_ _5141_/A _4965_/B vssd1 vssd1 vccd1 vccd1 _5118_/A sky130_fd_sc_hd__or2_1
XFILLER_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3916_ _7081_/A _5129_/A vssd1 vssd1 vccd1 vccd1 _3995_/B sky130_fd_sc_hd__nor2_1
X_6704_ _6960_/A _6704_/B _6704_/C vssd1 vssd1 vccd1 vccd1 _6704_/X sky130_fd_sc_hd__and3_1
XFILLER_51_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4896_ _4899_/A _4899_/B vssd1 vssd1 vccd1 vccd1 _4917_/B sky130_fd_sc_hd__nand2_1
XFILLER_32_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3847_ _7188_/Q _5674_/B vssd1 vssd1 vccd1 vccd1 _5267_/A sky130_fd_sc_hd__and2_2
X_6635_ _6635_/A _6635_/B vssd1 vssd1 vccd1 vccd1 _6636_/B sky130_fd_sc_hd__or2_1
X_6566_ _6566_/A _6566_/B vssd1 vssd1 vccd1 vccd1 _6568_/B sky130_fd_sc_hd__xnor2_2
X_3778_ _3778_/A vssd1 vssd1 vccd1 vccd1 _3783_/B sky130_fd_sc_hd__inv_2
X_5517_ _5560_/A _5560_/B vssd1 vssd1 vccd1 vccd1 _5520_/A sky130_fd_sc_hd__xnor2_1
X_6497_ _6487_/A _6487_/C _6487_/D _6487_/B vssd1 vssd1 vccd1 vccd1 _6497_/Y sky130_fd_sc_hd__a22oi_2
X_5448_ _5476_/A _5476_/B vssd1 vssd1 vccd1 vccd1 _5499_/A sky130_fd_sc_hd__xnor2_1
X_5379_ _5262_/X _5377_/X hold48/X _7226_/D vssd1 vssd1 vccd1 vccd1 hold49/A sky130_fd_sc_hd__o211a_1
XFILLER_101_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7118_ _7118_/A vssd1 vssd1 vccd1 vccd1 _7225_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7049_ _7025_/A _7045_/X _7047_/Y _7048_/X vssd1 vssd1 vccd1 vccd1 _7196_/D sky130_fd_sc_hd__o211a_1
XFILLER_27_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4750_ hold97/A _6687_/B _4593_/B _4679_/Y vssd1 vssd1 vccd1 vccd1 _4751_/B sky130_fd_sc_hd__o2bb2a_1
X_4681_ _4593_/B _4679_/Y hold97/A _4789_/B vssd1 vssd1 vccd1 vccd1 _4838_/B sky130_fd_sc_hd__and4bb_2
X_3701_ _3703_/A vssd1 vssd1 vccd1 vccd1 _3701_/Y sky130_fd_sc_hd__inv_2
X_3632_ _3635_/A vssd1 vssd1 vccd1 vccd1 _3632_/Y sky130_fd_sc_hd__inv_2
X_6420_ _6679_/A _6420_/B vssd1 vssd1 vccd1 vccd1 _6538_/A sky130_fd_sc_hd__nor2_1
X_6351_ _6351_/A _6351_/B vssd1 vssd1 vccd1 vccd1 _6352_/B sky130_fd_sc_hd__nor2_1
X_5302_ _7114_/A _6455_/A _5169_/Y vssd1 vssd1 vccd1 vccd1 _5304_/B sky130_fd_sc_hd__o21ai_1
XFILLER_88_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6282_ _6336_/A _6282_/B vssd1 vssd1 vccd1 vccd1 _6285_/A sky130_fd_sc_hd__xnor2_2
XFILLER_69_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5233_ _5015_/A _5015_/B _5006_/Y vssd1 vssd1 vccd1 vccd1 _5353_/B sky130_fd_sc_hd__o21ai_2
X_5164_ _5406_/A _6139_/A vssd1 vssd1 vccd1 vccd1 _5165_/B sky130_fd_sc_hd__nor2_1
X_4115_ _4115_/A _4230_/A vssd1 vssd1 vccd1 vccd1 _4117_/B sky130_fd_sc_hd__xnor2_1
XFILLER_83_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5095_ _5095_/A _5247_/B vssd1 vssd1 vccd1 vccd1 _5096_/B sky130_fd_sc_hd__xnor2_1
X_4046_ _7159_/Q vssd1 vssd1 vccd1 vccd1 _6016_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5997_ _5602_/A _5990_/Y _5996_/X _5990_/B vssd1 vssd1 vccd1 vccd1 _5998_/C sky130_fd_sc_hd__o211a_1
XFILLER_12_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4948_ _4948_/A _4948_/B vssd1 vssd1 vccd1 vccd1 _5111_/A sky130_fd_sc_hd__or2_2
X_4879_ _4891_/A _4891_/B vssd1 vssd1 vccd1 vccd1 _4892_/A sky130_fd_sc_hd__nand2_1
X_6618_ _6649_/A _6618_/B vssd1 vssd1 vccd1 vccd1 _6650_/A sky130_fd_sc_hd__nor2_1
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6549_ _6549_/A _6549_/B vssd1 vssd1 vccd1 vccd1 _6575_/B sky130_fd_sc_hd__xor2_2
X_7306__99 vssd1 vssd1 vccd1 vccd1 _7306__99/HI _7414_/A sky130_fd_sc_hd__conb_1
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5920_ _6994_/A _5918_/A _5948_/A _5944_/B _5919_/X vssd1 vssd1 vccd1 vccd1 _5924_/B
+ sky130_fd_sc_hd__o41ai_4
XFILLER_0_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5851_ _6162_/C vssd1 vssd1 vccd1 vccd1 _6301_/A sky130_fd_sc_hd__buf_2
X_4802_ _4802_/A _4802_/B _4802_/C vssd1 vssd1 vccd1 vccd1 _4819_/A sky130_fd_sc_hd__or3_2
X_5782_ _6537_/B _5782_/B vssd1 vssd1 vccd1 vccd1 _5789_/A sky130_fd_sc_hd__nand2_1
X_4733_ _4660_/Y _4733_/B vssd1 vssd1 vccd1 vccd1 _4734_/B sky130_fd_sc_hd__and2b_1
XFILLER_21_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4664_ _4686_/A _4686_/B vssd1 vssd1 vccd1 vccd1 _4689_/A sky130_fd_sc_hd__xnor2_1
X_6403_ _6403_/A _6403_/B vssd1 vssd1 vccd1 vccd1 _6403_/Y sky130_fd_sc_hd__nor2_1
X_3615_ _3616_/A vssd1 vssd1 vccd1 vccd1 _3615_/Y sky130_fd_sc_hd__inv_2
X_4595_ _4595_/A _4595_/B vssd1 vssd1 vccd1 vccd1 _4663_/B sky130_fd_sc_hd__xnor2_1
X_7383_ _7383_/A _3674_/Y vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_hd__ebufn_8
X_6334_ _7009_/A _7006_/A _7011_/A vssd1 vssd1 vccd1 vccd1 _6362_/B sky130_fd_sc_hd__o21a_1
XFILLER_88_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6265_ _6125_/A _6207_/B _6120_/A vssd1 vssd1 vccd1 vccd1 _6269_/A sky130_fd_sc_hd__a21o_1
XFILLER_88_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5216_ _5216_/A _5216_/B vssd1 vssd1 vccd1 vccd1 _5446_/B sky130_fd_sc_hd__nor2_1
X_6196_ _7117_/A vssd1 vssd1 vccd1 vccd1 _6196_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5147_ _5148_/A _5148_/B _5148_/C vssd1 vssd1 vccd1 vccd1 _5149_/A sky130_fd_sc_hd__a21oi_1
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5078_ _4147_/A _4147_/B _4150_/B vssd1 vssd1 vccd1 vccd1 _5236_/B sky130_fd_sc_hd__o21ai_2
X_4029_ _5131_/A _4193_/B _4028_/X vssd1 vssd1 vccd1 vccd1 _4189_/B sky130_fd_sc_hd__a21oi_2
XFILLER_25_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4380_ _4380_/A _5076_/A vssd1 vssd1 vccd1 vccd1 _4382_/C sky130_fd_sc_hd__xnor2_1
XFILLER_98_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6050_ _5710_/A _5710_/B _6049_/Y vssd1 vssd1 vccd1 vccd1 _6154_/B sky130_fd_sc_hd__a21oi_2
X_5001_ _3982_/A _5001_/B vssd1 vssd1 vccd1 vccd1 _5035_/B sky130_fd_sc_hd__and2b_1
XFILLER_66_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6952_ _7007_/A vssd1 vssd1 vccd1 vccd1 _6952_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5903_ _5991_/A _4796_/X _4328_/A _6241_/A vssd1 vssd1 vccd1 vccd1 _5938_/A sky130_fd_sc_hd__o211a_1
X_6883_ _6969_/A _6874_/B _6882_/X vssd1 vssd1 vccd1 vccd1 _6883_/Y sky130_fd_sc_hd__o21ai_1
X_5834_ _5871_/A _5832_/Y _5833_/Y vssd1 vssd1 vccd1 vccd1 _5835_/B sky130_fd_sc_hd__a21oi_1
XFILLER_34_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5765_ _5765_/A _6466_/B vssd1 vssd1 vccd1 vccd1 _5827_/B sky130_fd_sc_hd__xor2_2
X_4716_ _4717_/A _4717_/B vssd1 vssd1 vccd1 vccd1 _4936_/B sky130_fd_sc_hd__xor2_1
X_5696_ _5696_/A _5696_/B vssd1 vssd1 vccd1 vccd1 _5719_/B sky130_fd_sc_hd__xor2_4
X_4647_ _4857_/B _4542_/B _4646_/Y _4176_/B vssd1 vssd1 vccd1 vccd1 _4730_/B sky130_fd_sc_hd__o22a_1
X_7366_ _7366_/A _3652_/Y vssd1 vssd1 vccd1 vccd1 io_out[8] sky130_fd_sc_hd__ebufn_8
X_4578_ _4467_/B _4467_/C _5717_/A vssd1 vssd1 vccd1 vccd1 _4579_/B sky130_fd_sc_hd__a21oi_1
X_6317_ _6254_/B _6317_/B vssd1 vssd1 vccd1 vccd1 _6317_/X sky130_fd_sc_hd__and2b_1
X_6248_ _6182_/A _6182_/B _6247_/X vssd1 vssd1 vccd1 vccd1 _6314_/B sky130_fd_sc_hd__a21bo_1
X_6179_ _6180_/A _6180_/C _6180_/B vssd1 vssd1 vccd1 vccd1 _6250_/A sky130_fd_sc_hd__o21a_1
XFILLER_29_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 hold80/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold91 hold91/A vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_63_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3880_ _7214_/Q vssd1 vssd1 vccd1 vccd1 _5274_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5550_ _5551_/A _5551_/B _5551_/C vssd1 vssd1 vccd1 vccd1 _5552_/A sky130_fd_sc_hd__a21oi_1
X_4501_ _7185_/Q _7184_/Q vssd1 vssd1 vccd1 vccd1 _4613_/C sky130_fd_sc_hd__nor2_4
X_5481_ _5486_/B _5412_/C _5413_/B vssd1 vssd1 vccd1 vccd1 _5546_/A sky130_fd_sc_hd__o21ba_1
X_4432_ _6439_/B hold77/A vssd1 vssd1 vccd1 vccd1 _4659_/A sky130_fd_sc_hd__nor2b_2
X_7220_ _7221_/CLK _7220_/D vssd1 vssd1 vccd1 vccd1 _7220_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_0 _5190_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4363_ _4363_/A _4363_/B vssd1 vssd1 vccd1 vccd1 _5047_/B sky130_fd_sc_hd__xnor2_2
X_7151_ _7151_/CLK hold45/X vssd1 vssd1 vccd1 vccd1 _7390_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7082_ hold70/X _7075_/X _7081_/Y _7073_/X vssd1 vssd1 vccd1 vccd1 _7209_/D sky130_fd_sc_hd__o211a_1
X_4294_ _6722_/A _4226_/B _4293_/X vssd1 vssd1 vccd1 vccd1 _4303_/A sky130_fd_sc_hd__o21a_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6102_ _6102_/A _6102_/B vssd1 vssd1 vccd1 vccd1 _6102_/X sky130_fd_sc_hd__xor2_4
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6033_ _6033_/A _6033_/B vssd1 vssd1 vccd1 vccd1 _6129_/B sky130_fd_sc_hd__xnor2_2
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6935_ _6977_/A vssd1 vssd1 vccd1 vccd1 _6935_/X sky130_fd_sc_hd__clkbuf_2
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6866_ _6866_/A _6866_/B vssd1 vssd1 vccd1 vccd1 _6873_/B sky130_fd_sc_hd__and2_1
XFILLER_22_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6797_ _6797_/A _6797_/B _6797_/C vssd1 vssd1 vccd1 vccd1 _6799_/A sky130_fd_sc_hd__or3_1
X_5817_ _5643_/B _5603_/B _5614_/B _5636_/A _5801_/B vssd1 vssd1 vccd1 vccd1 _5818_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5748_ _5748_/A _5748_/B vssd1 vssd1 vccd1 vccd1 _6080_/B sky130_fd_sc_hd__xnor2_2
X_5679_ _5685_/A _5679_/B vssd1 vssd1 vccd1 vccd1 _6035_/B sky130_fd_sc_hd__xor2_2
X_7418_ _7418_/A _3711_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[22] sky130_fd_sc_hd__ebufn_8
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7349_ _7349_/A _3634_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[23] sky130_fd_sc_hd__ebufn_8
XFILLER_66_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4981_ _4981_/A _3891_/B vssd1 vssd1 vccd1 vccd1 _4992_/B sky130_fd_sc_hd__or2b_1
XFILLER_63_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3932_ _4019_/A _4019_/B _3931_/X vssd1 vssd1 vccd1 vccd1 _4996_/B sky130_fd_sc_hd__a21o_1
XFILLER_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6720_ _6720_/A _6720_/B vssd1 vssd1 vccd1 vccd1 _6722_/B sky130_fd_sc_hd__xnor2_1
X_3863_ _7196_/Q _7195_/Q vssd1 vssd1 vccd1 vccd1 _3998_/B sky130_fd_sc_hd__xor2_2
X_6651_ _6651_/A _6651_/B vssd1 vssd1 vccd1 vccd1 _6652_/A sky130_fd_sc_hd__nand2_1
XFILLER_31_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6582_ _6605_/A _6605_/B _6581_/X vssd1 vssd1 vccd1 vccd1 _6745_/A sky130_fd_sc_hd__a21oi_1
X_5602_ _5602_/A _5602_/B vssd1 vssd1 vccd1 vccd1 _5603_/B sky130_fd_sc_hd__or2_1
X_3794_ _4359_/B _3794_/B vssd1 vssd1 vccd1 vccd1 _4354_/A sky130_fd_sc_hd__xnor2_2
X_5533_ _5531_/X _5569_/B vssd1 vssd1 vccd1 vccd1 _5533_/X sky130_fd_sc_hd__and2b_1
X_5464_ _5464_/A _5464_/B vssd1 vssd1 vccd1 vccd1 _5464_/X sky130_fd_sc_hd__or2_1
X_4415_ _4416_/B _4415_/B vssd1 vssd1 vccd1 vccd1 _4538_/B sky130_fd_sc_hd__xnor2_1
X_7203_ _7222_/CLK _7203_/D vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__dfxtp_1
X_5395_ _5490_/A _5395_/B vssd1 vssd1 vccd1 vccd1 _5397_/C sky130_fd_sc_hd__nor2_1
X_7134_ _7224_/CLK _7134_/D vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__dfxtp_1
X_4346_ _7171_/Q vssd1 vssd1 vccd1 vccd1 _6563_/A sky130_fd_sc_hd__inv_2
XFILLER_101_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7065_ hold116/X _7062_/X _7064_/X _7060_/X vssd1 vssd1 vccd1 vccd1 _7202_/D sky130_fd_sc_hd__o211a_1
X_4277_ _4317_/A hold90/A vssd1 vssd1 vccd1 vccd1 _4278_/B sky130_fd_sc_hd__or2_1
X_6016_ _6016_/A _6439_/A vssd1 vssd1 vccd1 vccd1 _6266_/B sky130_fd_sc_hd__nand2_1
XFILLER_74_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7316__109 vssd1 vssd1 vccd1 vccd1 _7316__109/HI _7424_/A sky130_fd_sc_hd__conb_1
X_7281__74 vssd1 vssd1 vccd1 vccd1 _7281__74/HI _7380_/A sky130_fd_sc_hd__conb_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6918_ hold43/X _6893_/A _6917_/X vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__a21oi_1
XFILLER_42_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6849_ _6831_/A _6849_/B vssd1 vssd1 vccd1 vccd1 _6862_/A sky130_fd_sc_hd__and2b_1
XFILLER_52_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4200_ _4238_/A _4238_/B vssd1 vssd1 vccd1 vccd1 _4239_/A sky130_fd_sc_hd__or2_1
X_5180_ _5325_/A _5180_/B vssd1 vssd1 vccd1 vccd1 _5181_/B sky130_fd_sc_hd__xnor2_1
X_4131_ _5783_/B vssd1 vssd1 vccd1 vccd1 _5784_/B sky130_fd_sc_hd__clkbuf_2
X_4062_ _6494_/A vssd1 vssd1 vccd1 vccd1 _6938_/A sky130_fd_sc_hd__inv_2
XFILLER_36_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4964_ _4964_/A _4964_/B _4964_/C vssd1 vssd1 vccd1 vccd1 _4965_/B sky130_fd_sc_hd__nor3_1
X_3915_ _4412_/B vssd1 vssd1 vccd1 vccd1 _7081_/A sky130_fd_sc_hd__inv_2
X_6703_ _6686_/X _6700_/X _6702_/Y vssd1 vssd1 vccd1 vccd1 _6703_/X sky130_fd_sc_hd__o21ba_1
XFILLER_32_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4895_ _4895_/A _4895_/B _4895_/C _4895_/D vssd1 vssd1 vccd1 vccd1 _4899_/B sky130_fd_sc_hd__nand4_4
X_3846_ _7186_/Q _7185_/Q vssd1 vssd1 vccd1 vccd1 _3922_/B sky130_fd_sc_hd__xor2_4
X_6634_ _6665_/A _6634_/B vssd1 vssd1 vccd1 vccd1 _6635_/B sky130_fd_sc_hd__nor2_1
X_6565_ _6565_/A _6565_/B vssd1 vssd1 vccd1 vccd1 _6566_/B sky130_fd_sc_hd__xor2_1
X_3777_ _7173_/Q _7170_/Q vssd1 vssd1 vccd1 vccd1 _3778_/A sky130_fd_sc_hd__or2b_1
X_6496_ _6496_/A _6496_/B _6496_/C vssd1 vssd1 vccd1 vccd1 _6505_/A sky130_fd_sc_hd__or3_1
X_5516_ _5458_/A _5458_/B _5419_/A vssd1 vssd1 vccd1 vccd1 _5560_/B sky130_fd_sc_hd__a21oi_1
X_5447_ _5339_/A _5339_/B _5446_/X vssd1 vssd1 vccd1 vccd1 _5476_/B sky130_fd_sc_hd__o21ba_1
X_5378_ _5594_/A hold47/X vssd1 vssd1 vccd1 vccd1 hold48/A sky130_fd_sc_hd__or2_1
XFILLER_86_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7117_ _7117_/A _7117_/B vssd1 vssd1 vccd1 vccd1 _7118_/A sky130_fd_sc_hd__and2_1
X_4329_ _4329_/A _6613_/A vssd1 vssd1 vccd1 vccd1 _5854_/A sky130_fd_sc_hd__xnor2_4
X_7048_ _7073_/A vssd1 vssd1 vccd1 vccd1 _7048_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_101_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3700_ _3703_/A vssd1 vssd1 vccd1 vccd1 _3700_/Y sky130_fd_sc_hd__inv_2
X_4680_ hold98/X vssd1 vssd1 vccd1 vccd1 hold97/A sky130_fd_sc_hd__buf_2
X_3631_ _3635_/A vssd1 vssd1 vccd1 vccd1 _3631_/Y sky130_fd_sc_hd__inv_2
X_6350_ _6305_/A _6350_/B vssd1 vssd1 vccd1 vccd1 _6351_/B sky130_fd_sc_hd__and2b_1
X_5301_ _7114_/A _6174_/A _5287_/A _5173_/B vssd1 vssd1 vccd1 vccd1 _5307_/A sky130_fd_sc_hd__o31a_1
X_6281_ _7011_/A _6141_/X _7006_/A vssd1 vssd1 vccd1 vccd1 _6282_/B sky130_fd_sc_hd__mux2_1
X_5232_ _6129_/A _5232_/B vssd1 vssd1 vccd1 vccd1 _5234_/A sky130_fd_sc_hd__xnor2_1
X_5163_ _5690_/A _5719_/A vssd1 vssd1 vccd1 vccd1 _6139_/A sky130_fd_sc_hd__and2_1
XFILLER_96_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4114_ _4317_/A _7167_/Q vssd1 vssd1 vccd1 vccd1 _4230_/A sky130_fd_sc_hd__nand2_1
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5094_ _5246_/B _5094_/B vssd1 vssd1 vccd1 vccd1 _5247_/B sky130_fd_sc_hd__xnor2_1
XFILLER_83_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4045_ _4045_/A _5039_/A vssd1 vssd1 vccd1 vccd1 _4167_/A sky130_fd_sc_hd__xnor2_2
XFILLER_37_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7251__44 vssd1 vssd1 vccd1 vccd1 _7251__44/HI _7350_/A sky130_fd_sc_hd__conb_1
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5996_ _5602_/A _5990_/Y _5995_/Y _5989_/B vssd1 vssd1 vccd1 vccd1 _5996_/X sky130_fd_sc_hd__a211o_1
XFILLER_52_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4947_ _3750_/X hold15/X _3752_/X _4946_/X vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__o211a_1
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4878_ _4878_/A _4878_/B vssd1 vssd1 vccd1 vccd1 _4891_/B sky130_fd_sc_hd__and2_1
XFILLER_20_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3829_ _5145_/A _5145_/B vssd1 vssd1 vccd1 vccd1 _3832_/B sky130_fd_sc_hd__xnor2_1
X_6617_ _6617_/A _6651_/A vssd1 vssd1 vccd1 vccd1 _6618_/B sky130_fd_sc_hd__and2_1
X_6548_ _6571_/A _6571_/B _6547_/A vssd1 vssd1 vccd1 vccd1 _6549_/B sky130_fd_sc_hd__a21o_1
X_6479_ _6588_/A _6479_/B vssd1 vssd1 vccd1 vccd1 _6480_/C sky130_fd_sc_hd__nor2_1
XFILLER_58_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5850_ _6409_/A _5850_/B vssd1 vssd1 vccd1 vccd1 _5857_/A sky130_fd_sc_hd__nand2_1
X_4801_ _4728_/B _4728_/C hold71/A vssd1 vssd1 vccd1 vccd1 _4802_/C sky130_fd_sc_hd__a21oi_1
X_5781_ _5758_/A _5838_/B _5755_/B vssd1 vssd1 vccd1 vccd1 _6085_/B sky130_fd_sc_hd__o21ai_2
X_4732_ _4770_/A _4770_/B vssd1 vssd1 vccd1 vccd1 _4771_/A sky130_fd_sc_hd__nor2_1
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4663_ _4663_/A _4663_/B vssd1 vssd1 vccd1 vccd1 _4686_/B sky130_fd_sc_hd__xor2_1
X_3614_ _3616_/A vssd1 vssd1 vccd1 vccd1 _3614_/Y sky130_fd_sc_hd__inv_2
X_6402_ _6402_/A _6402_/B vssd1 vssd1 vccd1 vccd1 _6403_/B sky130_fd_sc_hd__xnor2_1
X_4594_ hold91/A _6620_/A _4785_/B vssd1 vssd1 vccd1 vccd1 _4595_/B sky130_fd_sc_hd__a21oi_1
X_7382_ _7382_/A _3672_/Y vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__ebufn_8
X_6333_ _6365_/A _6333_/B vssd1 vssd1 vccd1 vccd1 _6335_/A sky130_fd_sc_hd__or2_1
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6264_ _6264_/A _6264_/B vssd1 vssd1 vccd1 vccd1 _6274_/B sky130_fd_sc_hd__nand2_1
X_5215_ _5215_/A _5215_/B _5215_/C vssd1 vssd1 vccd1 vccd1 _5216_/B sky130_fd_sc_hd__and3_1
X_6195_ _6391_/A hold37/X vssd1 vssd1 vccd1 vccd1 _6195_/X sky130_fd_sc_hd__or2_1
X_5146_ _5287_/A _5146_/B vssd1 vssd1 vccd1 vccd1 _5148_/C sky130_fd_sc_hd__xnor2_1
XFILLER_29_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5077_ _5229_/A _4379_/B _5076_/X vssd1 vssd1 vccd1 vccd1 _5088_/A sky130_fd_sc_hd__o21ai_2
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4028_ _4426_/A _7211_/Q vssd1 vssd1 vccd1 vccd1 _4028_/X sky130_fd_sc_hd__and2_1
XFILLER_25_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5979_ _5978_/A _5986_/A _5983_/B _5983_/A vssd1 vssd1 vccd1 vccd1 _5980_/B sky130_fd_sc_hd__o22a_1
XFILLER_40_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5000_ _3981_/B _5000_/B vssd1 vssd1 vccd1 vccd1 _5035_/A sky130_fd_sc_hd__and2b_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6951_ _7020_/A vssd1 vssd1 vccd1 vccd1 _7007_/A sky130_fd_sc_hd__clkbuf_2
X_5902_ _5915_/A _5902_/B vssd1 vssd1 vccd1 vccd1 _5922_/A sky130_fd_sc_hd__xnor2_1
X_6882_ _6969_/A _6874_/B _6875_/A _6875_/B vssd1 vssd1 vccd1 vccd1 _6882_/X sky130_fd_sc_hd__a22o_1
X_5833_ _5833_/A _5833_/B vssd1 vssd1 vccd1 vccd1 _5833_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5764_ _6502_/A vssd1 vssd1 vccd1 vccd1 _6466_/B sky130_fd_sc_hd__clkbuf_2
X_4715_ _4720_/A _4720_/B _4714_/Y vssd1 vssd1 vccd1 vccd1 _4717_/B sky130_fd_sc_hd__a21oi_1
X_5695_ _5696_/A _5696_/B vssd1 vssd1 vccd1 vccd1 _5698_/A sky130_fd_sc_hd__nand2_1
XFILLER_30_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4646_ _4799_/B _4726_/B vssd1 vssd1 vccd1 vccd1 _4646_/Y sky130_fd_sc_hd__nor2_1
X_4577_ _5827_/A vssd1 vssd1 vccd1 vccd1 _5717_/A sky130_fd_sc_hd__buf_2
XFILLER_30_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7365_ _7365_/A _3651_/Y vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__ebufn_8
XFILLER_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6316_ _6316_/A _6357_/B vssd1 vssd1 vccd1 vccd1 _6319_/A sky130_fd_sc_hd__xnor2_2
X_6247_ _6247_/A _6173_/A vssd1 vssd1 vccd1 vccd1 _6247_/X sky130_fd_sc_hd__or2b_1
XFILLER_39_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6178_ _6075_/A _6074_/A _6167_/B _6078_/B vssd1 vssd1 vccd1 vccd1 _6180_/B sky130_fd_sc_hd__a31o_1
XFILLER_84_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5129_ _5129_/A vssd1 vssd1 vccd1 vccd1 _5478_/A sky130_fd_sc_hd__buf_2
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7287__80 vssd1 vssd1 vccd1 vccd1 _7287__80/HI _7395_/A sky130_fd_sc_hd__conb_1
XFILLER_88_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold92 hold92/A vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold70/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_75_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4500_ _4500_/A _4500_/B vssd1 vssd1 vccd1 vccd1 _4511_/A sky130_fd_sc_hd__xnor2_2
X_5480_ _6240_/A _5168_/X _5143_/X _7114_/A vssd1 vssd1 vccd1 vccd1 _5486_/B sky130_fd_sc_hd__o2bb2a_1
XANTENNA_1 _4520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4431_ _5691_/B vssd1 vssd1 vccd1 vccd1 _6439_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4362_ _5055_/A _5056_/D vssd1 vssd1 vccd1 vccd1 _4363_/B sky130_fd_sc_hd__xor2_1
X_7150_ _7151_/CLK hold7/X vssd1 vssd1 vccd1 vccd1 _7389_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_98_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7081_ _7081_/A _7093_/B vssd1 vssd1 vccd1 vccd1 _7081_/Y sky130_fd_sc_hd__nand2_1
XFILLER_86_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4293_ _4293_/A _4233_/B vssd1 vssd1 vccd1 vccd1 _4293_/X sky130_fd_sc_hd__or2b_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6101_ _6011_/A _6011_/B _6100_/X vssd1 vssd1 vccd1 vccd1 _6102_/B sky130_fd_sc_hd__a21o_2
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6032_ _6128_/B _6116_/B vssd1 vssd1 vccd1 vccd1 _6033_/B sky130_fd_sc_hd__xnor2_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6934_ input4/X _7116_/B _6933_/Y _6846_/X vssd1 vssd1 vccd1 vccd1 _7155_/D sky130_fd_sc_hd__o211a_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6865_ _6865_/A _6836_/B vssd1 vssd1 vccd1 vccd1 _6866_/B sky130_fd_sc_hd__or2b_1
X_6796_ _6796_/A _6796_/B vssd1 vssd1 vccd1 vccd1 _6797_/C sky130_fd_sc_hd__xnor2_1
X_5816_ _5849_/B _5816_/B vssd1 vssd1 vccd1 vccd1 _5819_/B sky130_fd_sc_hd__xor2_1
XFILLER_22_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5747_ _5747_/A _5747_/B vssd1 vssd1 vccd1 vccd1 _5748_/B sky130_fd_sc_hd__and2_1
X_7417_ _7417_/A _3713_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[21] sky130_fd_sc_hd__ebufn_8
X_5678_ _6029_/B _5678_/B vssd1 vssd1 vccd1 vccd1 _5679_/B sky130_fd_sc_hd__xor2_2
X_4629_ _4629_/A _4629_/B vssd1 vssd1 vccd1 vccd1 _4629_/Y sky130_fd_sc_hd__nor2_1
X_7348_ _7348_/A _3633_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[22] sky130_fd_sc_hd__ebufn_8
XFILLER_89_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4980_ _3980_/A _3980_/B _3979_/A vssd1 vssd1 vccd1 vccd1 _4994_/A sky130_fd_sc_hd__a21o_1
XFILLER_16_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3931_ _3931_/A _3931_/B vssd1 vssd1 vccd1 vccd1 _3931_/X sky130_fd_sc_hd__and2_1
X_3862_ _7197_/Q vssd1 vssd1 vccd1 vccd1 _3910_/A sky130_fd_sc_hd__clkbuf_2
X_6650_ _6650_/A _6650_/B vssd1 vssd1 vccd1 vccd1 _6706_/C sky130_fd_sc_hd__xnor2_1
X_6581_ _6580_/B _6581_/B vssd1 vssd1 vccd1 vccd1 _6581_/X sky130_fd_sc_hd__and2b_1
X_5601_ _5602_/A _5602_/B vssd1 vssd1 vccd1 vccd1 _5643_/B sky130_fd_sc_hd__nand2_2
X_3793_ _7066_/A _4356_/B _4359_/A vssd1 vssd1 vccd1 vccd1 _3794_/B sky130_fd_sc_hd__o21ai_1
X_5532_ _5531_/A _5531_/B _5531_/C vssd1 vssd1 vccd1 vccd1 _5569_/B sky130_fd_sc_hd__a21o_1
X_5463_ _5463_/A _5463_/B vssd1 vssd1 vccd1 vccd1 _5466_/A sky130_fd_sc_hd__xor2_1
XFILLER_99_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4414_ _3879_/B _4649_/B _4413_/X vssd1 vssd1 vccd1 vccd1 _4415_/B sky130_fd_sc_hd__o21a_1
X_7202_ _7221_/CLK _7202_/D vssd1 vssd1 vccd1 vccd1 _7202_/Q sky130_fd_sc_hd__dfxtp_1
X_5394_ _5394_/A _5394_/B _5394_/C vssd1 vssd1 vccd1 vccd1 _5395_/B sky130_fd_sc_hd__and3_1
X_7133_ _7224_/CLK _7133_/D vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfxtp_1
X_4345_ _4477_/A vssd1 vssd1 vccd1 vccd1 _5218_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4276_ _4310_/A vssd1 vssd1 vccd1 vccd1 _5812_/A sky130_fd_sc_hd__buf_2
X_7064_ hold91/X _7091_/B vssd1 vssd1 vccd1 vccd1 _7064_/X sky130_fd_sc_hd__or2_1
XFILLER_59_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6015_ _5682_/A _5682_/B _5664_/B _6014_/Y vssd1 vssd1 vccd1 vccd1 _6107_/A sky130_fd_sc_hd__a31oi_4
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6917_ hold14/X _6893_/B _6894_/A hold23/X vssd1 vssd1 vccd1 vccd1 _6917_/X sky130_fd_sc_hd__a22o_1
X_6848_ _6839_/A _6848_/B vssd1 vssd1 vccd1 vccd1 _6869_/A sky130_fd_sc_hd__and2b_1
XFILLER_50_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6779_ _6744_/A _6778_/Y _6743_/A vssd1 vssd1 vccd1 vccd1 _6792_/B sky130_fd_sc_hd__o21a_1
XFILLER_2_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7257__50 vssd1 vssd1 vccd1 vccd1 _7257__50/HI _7356_/A sky130_fd_sc_hd__conb_1
XFILLER_77_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4130_ _7167_/Q vssd1 vssd1 vccd1 vccd1 _5783_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4061_ _5017_/A _4152_/C vssd1 vssd1 vccd1 vccd1 _4064_/A sky130_fd_sc_hd__nor2_1
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4963_ _4964_/A _4964_/B _4964_/C vssd1 vssd1 vccd1 vccd1 _5141_/A sky130_fd_sc_hd__o21a_1
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3914_ _4412_/B _4956_/B vssd1 vssd1 vccd1 vccd1 _3995_/A sky130_fd_sc_hd__and2b_1
X_6702_ _6686_/X _6700_/X _6701_/X vssd1 vssd1 vccd1 vccd1 _6702_/Y sky130_fd_sc_hd__a21oi_1
X_4894_ _7036_/A _7014_/A vssd1 vssd1 vccd1 vccd1 _4895_/D sky130_fd_sc_hd__or2_1
X_6633_ _6631_/A _6631_/B _6654_/A vssd1 vssd1 vccd1 vccd1 _6637_/B sky130_fd_sc_hd__o21ai_2
XFILLER_20_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3845_ _4011_/A _4011_/B _3844_/X vssd1 vssd1 vccd1 vccd1 _4252_/A sky130_fd_sc_hd__o21ai_4
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6564_ _6564_/A vssd1 vssd1 vccd1 vccd1 _6981_/A sky130_fd_sc_hd__clkinv_2
X_3776_ _5615_/A _5625_/A vssd1 vssd1 vccd1 vccd1 _3783_/A sky130_fd_sc_hd__nor2_1
X_6495_ _6502_/A _6502_/B _6483_/A vssd1 vssd1 vccd1 vccd1 _6496_/C sky130_fd_sc_hd__a21oi_1
X_5515_ _5515_/A _5537_/B vssd1 vssd1 vccd1 vccd1 _5560_/A sky130_fd_sc_hd__xor2_1
X_5446_ _5446_/A _5446_/B _5446_/C vssd1 vssd1 vccd1 vccd1 _5446_/X sky130_fd_sc_hd__and3_1
XFILLER_87_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5377_ _5375_/X _5472_/B vssd1 vssd1 vccd1 vccd1 _5377_/X sky130_fd_sc_hd__and2b_1
X_4328_ _4328_/A _4328_/B vssd1 vssd1 vccd1 vccd1 _4330_/A sky130_fd_sc_hd__nand2_1
X_7116_ _7116_/A _7116_/B vssd1 vssd1 vccd1 vccd1 _7224_/D sky130_fd_sc_hd__nor2_1
X_7047_ _7047_/A _7072_/B vssd1 vssd1 vccd1 vccd1 _7047_/Y sky130_fd_sc_hd__nand2_1
XFILLER_101_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4259_ _4259_/A _4260_/C vssd1 vssd1 vccd1 vccd1 _4494_/B sky130_fd_sc_hd__xnor2_2
XFILLER_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3630_ _3648_/A vssd1 vssd1 vccd1 vccd1 _3635_/A sky130_fd_sc_hd__clkbuf_16
X_5300_ _5611_/C vssd1 vssd1 vccd1 vccd1 _6174_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6280_ _6280_/A _6280_/B vssd1 vssd1 vccd1 vccd1 _6336_/A sky130_fd_sc_hd__xnor2_2
X_5231_ _5231_/A _5231_/B vssd1 vssd1 vccd1 vccd1 _5232_/B sky130_fd_sc_hd__nor2_1
X_5162_ _5689_/A _6140_/A _5784_/B vssd1 vssd1 vccd1 vccd1 _5348_/S sky130_fd_sc_hd__and3_1
XFILLER_68_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5093_ _5093_/A _5093_/B vssd1 vssd1 vccd1 vccd1 _5094_/B sky130_fd_sc_hd__xnor2_1
X_4113_ _7179_/Q vssd1 vssd1 vccd1 vccd1 _4317_/A sky130_fd_sc_hd__buf_4
X_4044_ _4044_/A _4044_/B vssd1 vssd1 vccd1 vccd1 _5039_/A sky130_fd_sc_hd__nor2_1
XFILLER_83_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5995_ _6950_/A _5987_/C _5994_/X vssd1 vssd1 vccd1 vccd1 _5995_/Y sky130_fd_sc_hd__o21ai_1
X_4946_ _4942_/Y _5111_/B hold63/X vssd1 vssd1 vccd1 vccd1 _4946_/X sky130_fd_sc_hd__a21o_1
X_4877_ _4858_/A _4858_/B _4895_/A vssd1 vssd1 vccd1 vccd1 _4878_/B sky130_fd_sc_hd__o21ai_1
X_3828_ _7089_/A _5273_/A _3827_/Y vssd1 vssd1 vccd1 vccd1 _5145_/B sky130_fd_sc_hd__o21a_1
XFILLER_20_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6616_ _6617_/A _6651_/A vssd1 vssd1 vccd1 vccd1 _6649_/A sky130_fd_sc_hd__nor2_1
X_6547_ _6547_/A _6547_/B vssd1 vssd1 vccd1 vccd1 _6571_/B sky130_fd_sc_hd__nor2_1
X_3759_ _7172_/Q vssd1 vssd1 vccd1 vccd1 _5198_/B sky130_fd_sc_hd__clkbuf_2
X_6478_ _6765_/A _6765_/B _6766_/A vssd1 vssd1 vccd1 vccd1 _6797_/A sky130_fd_sc_hd__a21boi_2
XFILLER_79_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5429_ _5784_/A _5430_/A vssd1 vssd1 vccd1 vccd1 _5432_/A sky130_fd_sc_hd__or2_1
XFILLER_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7227__20 vssd1 vssd1 vccd1 vccd1 _7227__20/HI _7326_/A sky130_fd_sc_hd__conb_1
XFILLER_74_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4800_ _4856_/A _4856_/B vssd1 vssd1 vccd1 vccd1 _4802_/B sky130_fd_sc_hd__nand2_1
XFILLER_21_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5780_ _6080_/B _5780_/B vssd1 vssd1 vccd1 vccd1 _5811_/A sky130_fd_sc_hd__xnor2_2
X_4731_ _4731_/A _4731_/B vssd1 vssd1 vccd1 vccd1 _4770_/B sky130_fd_sc_hd__or2_1
XFILLER_14_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4662_ _4691_/A _4734_/A _4656_/A vssd1 vssd1 vccd1 vccd1 _4686_/A sky130_fd_sc_hd__a21o_1
X_3613_ _3616_/A vssd1 vssd1 vccd1 vccd1 _3613_/Y sky130_fd_sc_hd__inv_2
X_6401_ _6401_/A _6401_/B vssd1 vssd1 vccd1 vccd1 _6402_/B sky130_fd_sc_hd__xnor2_1
X_4593_ _4838_/A _4593_/B vssd1 vssd1 vccd1 vccd1 _4785_/B sky130_fd_sc_hd__and2_1
X_7381_ _7381_/A _3671_/Y vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__ebufn_8
X_6332_ _6332_/A _6332_/B _6332_/C vssd1 vssd1 vccd1 vccd1 _6333_/B sky130_fd_sc_hd__nor3_1
X_6263_ _6263_/A _6263_/B vssd1 vssd1 vccd1 vccd1 _6274_/A sky130_fd_sc_hd__nand2_1
X_5214_ _5215_/A _5215_/B _5215_/C vssd1 vssd1 vccd1 vccd1 _5216_/A sky130_fd_sc_hd__a21oi_1
X_6194_ _6194_/A _6194_/B vssd1 vssd1 vccd1 vccd1 _6194_/X sky130_fd_sc_hd__xor2_4
XFILLER_84_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5145_ _5145_/A _5145_/B _5145_/C vssd1 vssd1 vccd1 vccd1 _5148_/A sky130_fd_sc_hd__or3_1
XFILLER_56_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5076_ _5076_/A _4380_/A vssd1 vssd1 vccd1 vccd1 _5076_/X sky130_fd_sc_hd__or2b_1
X_4027_ _4426_/A _7211_/Q vssd1 vssd1 vccd1 vccd1 _4193_/B sky130_fd_sc_hd__xor2_2
XFILLER_71_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5978_ _5978_/A _5978_/B vssd1 vssd1 vccd1 vccd1 _5983_/B sky130_fd_sc_hd__xor2_1
X_4929_ _4932_/A _4932_/B vssd1 vssd1 vccd1 vccd1 _4929_/Y sky130_fd_sc_hd__nand2_1
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6950_ _6950_/A _6954_/B vssd1 vssd1 vccd1 vccd1 _6950_/X sky130_fd_sc_hd__or2_1
XFILLER_81_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5901_ _5914_/A _5914_/B vssd1 vssd1 vccd1 vccd1 _5915_/A sky130_fd_sc_hd__nor2_1
XFILLER_53_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6881_ _6906_/A hold66/X vssd1 vssd1 vccd1 vccd1 _7142_/D sky130_fd_sc_hd__nor2_1
XFILLER_34_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5832_ _5871_/B vssd1 vssd1 vccd1 vccd1 _5832_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5763_ _7154_/Q vssd1 vssd1 vccd1 vccd1 _6502_/A sky130_fd_sc_hd__clkbuf_2
X_4714_ _4714_/A _4714_/B vssd1 vssd1 vccd1 vccd1 _4714_/Y sky130_fd_sc_hd__nor2_1
X_5694_ _5694_/A _5723_/A vssd1 vssd1 vccd1 vccd1 _5696_/B sky130_fd_sc_hd__xnor2_4
X_4645_ _4659_/B _4645_/B vssd1 vssd1 vccd1 vccd1 _4730_/A sky130_fd_sc_hd__nor2_1
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7433_ _7433_/A _3732_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[37] sky130_fd_sc_hd__ebufn_8
X_7364_ _7364_/A _3650_/Y vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__ebufn_8
X_4576_ _4914_/B _4668_/B vssd1 vssd1 vccd1 vccd1 _4580_/A sky130_fd_sc_hd__nand2_1
X_6315_ _6250_/A _6250_/B _6314_/Y vssd1 vssd1 vccd1 vccd1 _6357_/B sky130_fd_sc_hd__a21bo_1
XFILLER_89_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6246_ _6246_/A _6246_/B vssd1 vssd1 vccd1 vccd1 _6314_/A sky130_fd_sc_hd__xnor2_1
X_6177_ _6177_/A _6245_/A vssd1 vssd1 vccd1 vccd1 _6180_/C sky130_fd_sc_hd__and2_1
XFILLER_84_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5128_ _5284_/A _5128_/B vssd1 vssd1 vccd1 vccd1 _5266_/A sky130_fd_sc_hd__nor2_1
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5059_ hold83/A hold87/A vssd1 vssd1 vccd1 vccd1 _5209_/B sky130_fd_sc_hd__xor2_1
XFILLER_55_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold71/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold82 hold82/A vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_90_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_90_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4430_ _7152_/Q vssd1 vssd1 vccd1 vccd1 _5691_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA_2 _6620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4361_ _5062_/C _4361_/B vssd1 vssd1 vccd1 vccd1 _5056_/D sky130_fd_sc_hd__xnor2_1
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6100_ _5934_/A _6100_/B vssd1 vssd1 vccd1 vccd1 _6100_/X sky130_fd_sc_hd__and2b_1
X_7080_ _7080_/A vssd1 vssd1 vccd1 vccd1 _7093_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4292_ _4334_/A _4334_/B _4291_/X vssd1 vssd1 vccd1 vccd1 _4304_/A sky130_fd_sc_hd__a21o_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6031_ _6118_/B _6031_/B vssd1 vssd1 vccd1 vccd1 _6116_/B sky130_fd_sc_hd__xnor2_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6933_ _6933_/A _6933_/B vssd1 vssd1 vccd1 vccd1 _6933_/Y sky130_fd_sc_hd__nand2_1
XFILLER_54_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6864_ _6864_/A _6835_/A vssd1 vssd1 vccd1 vccd1 _6866_/A sky130_fd_sc_hd__or2b_1
XFILLER_34_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5815_ _5815_/A _5815_/B vssd1 vssd1 vccd1 vccd1 _5816_/B sky130_fd_sc_hd__xnor2_2
X_6795_ _6758_/B _6761_/Y _6865_/A vssd1 vssd1 vccd1 vccd1 _6808_/A sky130_fd_sc_hd__o21a_1
X_5746_ _5745_/A _5745_/B _5745_/C vssd1 vssd1 vccd1 vccd1 _5747_/B sky130_fd_sc_hd__o21ai_1
X_5677_ _5669_/B _5669_/C _6029_/A vssd1 vssd1 vccd1 vccd1 _5678_/B sky130_fd_sc_hd__o21a_1
X_4628_ _4629_/A _4629_/B vssd1 vssd1 vccd1 vccd1 _4636_/B sky130_fd_sc_hd__xor2_1
X_7416_ _7416_/A _3715_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[20] sky130_fd_sc_hd__ebufn_8
X_4559_ _4559_/A _4559_/B vssd1 vssd1 vccd1 vccd1 _4560_/B sky130_fd_sc_hd__xor2_1
X_7347_ _7347_/A _3632_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[21] sky130_fd_sc_hd__ebufn_8
X_6229_ _6420_/B _6228_/C _6962_/A vssd1 vssd1 vccd1 vccd1 _6230_/B sky130_fd_sc_hd__a21oi_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3930_ _3931_/A _3931_/B vssd1 vssd1 vccd1 vccd1 _4019_/B sky130_fd_sc_hd__xor2_2
XFILLER_16_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3861_ _4956_/B _3861_/B vssd1 vssd1 vccd1 vccd1 _3867_/A sky130_fd_sc_hd__xnor2_1
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3792_ _7201_/Q _7204_/Q vssd1 vssd1 vccd1 vccd1 _4359_/A sky130_fd_sc_hd__or2b_1
X_6580_ _6581_/B _6580_/B vssd1 vssd1 vccd1 vccd1 _6605_/B sky130_fd_sc_hd__xnor2_1
X_5600_ _5804_/A _5796_/B _5640_/A vssd1 vssd1 vccd1 vccd1 _5602_/B sky130_fd_sc_hd__mux2_1
X_5531_ _5531_/A _5531_/B _5531_/C vssd1 vssd1 vccd1 vccd1 _5531_/X sky130_fd_sc_hd__and3_1
X_7201_ _7222_/CLK _7201_/D vssd1 vssd1 vccd1 vccd1 _7201_/Q sky130_fd_sc_hd__dfxtp_1
X_5462_ _5358_/A _5358_/B _5461_/X vssd1 vssd1 vccd1 vccd1 _5463_/B sky130_fd_sc_hd__a21boi_1
X_4413_ _7085_/A _4540_/B _4541_/B vssd1 vssd1 vccd1 vccd1 _4413_/X sky130_fd_sc_hd__or3_1
X_5393_ _5394_/A _5394_/B _5394_/C vssd1 vssd1 vccd1 vccd1 _5490_/A sky130_fd_sc_hd__a21oi_2
X_7132_ _7224_/CLK _7132_/D vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__dfxtp_1
X_4344_ _4344_/A _4344_/B vssd1 vssd1 vccd1 vccd1 _4366_/A sky130_fd_sc_hd__nor2_2
XFILLER_98_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7063_ _7063_/A vssd1 vssd1 vccd1 vccd1 _7091_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6014_ _6014_/A _6014_/B _6020_/B vssd1 vssd1 vccd1 vccd1 _6014_/Y sky130_fd_sc_hd__nor3_1
X_4275_ hold90/A _5734_/A vssd1 vssd1 vccd1 vccd1 _4310_/A sky130_fd_sc_hd__nand2_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6916_ _7116_/A hold8/X vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__nor2_1
XFILLER_35_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6847_ _6261_/X _6844_/Y hold67/X _6846_/X vssd1 vssd1 vccd1 vccd1 hold69/A sky130_fd_sc_hd__o211a_1
XFILLER_52_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6778_ _6778_/A _6778_/B _6778_/C vssd1 vssd1 vccd1 vccd1 _6778_/Y sky130_fd_sc_hd__nor3_1
XFILLER_22_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5729_ _5760_/A _5760_/B _5728_/X vssd1 vssd1 vccd1 vccd1 _5730_/B sky130_fd_sc_hd__o21ba_2
XFILLER_22_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7272__65 vssd1 vssd1 vccd1 vccd1 _7272__65/HI _7371_/A sky130_fd_sc_hd__conb_1
XFILLER_18_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4060_ _5597_/B _6449_/A vssd1 vssd1 vccd1 vccd1 _4152_/C sky130_fd_sc_hd__and2_1
XFILLER_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4962_ _5119_/A _5120_/B vssd1 vssd1 vccd1 vccd1 _4964_/C sky130_fd_sc_hd__xnor2_1
X_3913_ _7209_/Q vssd1 vssd1 vccd1 vccd1 _4412_/B sky130_fd_sc_hd__clkbuf_2
X_4893_ hold80/A _7078_/A vssd1 vssd1 vccd1 vccd1 _4895_/C sky130_fd_sc_hd__or2_1
X_6701_ _6701_/A _6701_/B vssd1 vssd1 vccd1 vccd1 _6701_/X sky130_fd_sc_hd__xor2_1
X_3844_ _4009_/A vssd1 vssd1 vccd1 vccd1 _3844_/X sky130_fd_sc_hd__clkbuf_2
X_6632_ _6947_/A _6653_/B vssd1 vssd1 vccd1 vccd1 _6654_/A sky130_fd_sc_hd__or2_1
XFILLER_20_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6563_ _6563_/A vssd1 vssd1 vccd1 vccd1 _6978_/A sky130_fd_sc_hd__buf_2
X_3775_ _7170_/Q vssd1 vssd1 vccd1 vccd1 _5625_/A sky130_fd_sc_hd__clkbuf_2
X_6494_ _6494_/A _6494_/B _7153_/Q vssd1 vssd1 vccd1 vccd1 _6496_/A sky130_fd_sc_hd__and3_1
X_5514_ _5558_/B _5514_/B vssd1 vssd1 vccd1 vccd1 _5537_/B sky130_fd_sc_hd__and2_1
X_7322__115 vssd1 vssd1 vccd1 vccd1 _7322__115/HI _7430_/A sky130_fd_sc_hd__conb_1
X_5445_ _5575_/A _5445_/B vssd1 vssd1 vccd1 vccd1 _5476_/A sky130_fd_sc_hd__nand2_1
X_7115_ _7096_/A _6933_/B _7114_/X _6405_/X vssd1 vssd1 vccd1 vccd1 _7223_/D sky130_fd_sc_hd__o211a_1
X_5376_ _5375_/A _5375_/B _5375_/C vssd1 vssd1 vccd1 vccd1 _5472_/B sky130_fd_sc_hd__a21o_1
XFILLER_87_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4327_ _4794_/A _4573_/A vssd1 vssd1 vccd1 vccd1 _4328_/B sky130_fd_sc_hd__or2_2
X_4258_ _4497_/A _4497_/B _4257_/X vssd1 vssd1 vccd1 vccd1 _4260_/C sky130_fd_sc_hd__o21a_1
X_7046_ _7080_/A vssd1 vssd1 vccd1 vccd1 _7072_/B sky130_fd_sc_hd__clkbuf_2
X_4189_ _4189_/A _4189_/B vssd1 vssd1 vccd1 vccd1 _4195_/A sky130_fd_sc_hd__xnor2_2
XFILLER_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5230_ _5229_/B _5229_/C _5229_/A vssd1 vssd1 vccd1 vccd1 _5231_/B sky130_fd_sc_hd__a21oi_1
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5161_ _5161_/A vssd1 vssd1 vccd1 vccd1 _6850_/A sky130_fd_sc_hd__buf_4
XFILLER_96_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5092_ _5092_/A _5092_/B vssd1 vssd1 vccd1 vccd1 _5093_/B sky130_fd_sc_hd__nor2_1
X_4112_ _6713_/A _4377_/B vssd1 vssd1 vccd1 vccd1 _4115_/A sky130_fd_sc_hd__xnor2_1
X_4043_ _4237_/A _4237_/B vssd1 vssd1 vccd1 vccd1 _4044_/B sky130_fd_sc_hd__and2b_1
XFILLER_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5994_ _5987_/A _6971_/A _5991_/A _5987_/C _5993_/X vssd1 vssd1 vccd1 vccd1 _5994_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_37_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4945_ hold74/X vssd1 vssd1 vccd1 vccd1 hold63/A sky130_fd_sc_hd__clkbuf_4
XFILLER_24_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4876_ _4876_/A _4895_/B vssd1 vssd1 vccd1 vccd1 _4891_/A sky130_fd_sc_hd__xor2_1
X_3827_ _4527_/A _3851_/B vssd1 vssd1 vccd1 vccd1 _3827_/Y sky130_fd_sc_hd__nand2_1
X_6615_ _6619_/A _6619_/B vssd1 vssd1 vccd1 vccd1 _6651_/A sky130_fd_sc_hd__or2_2
X_3758_ _7172_/Q _5625_/B vssd1 vssd1 vccd1 vccd1 _3761_/B sky130_fd_sc_hd__or2_1
X_6546_ _6546_/A _6546_/B vssd1 vssd1 vccd1 vccd1 _6547_/B sky130_fd_sc_hd__nor2_1
X_3689_ _3691_/A vssd1 vssd1 vccd1 vccd1 _3689_/Y sky130_fd_sc_hd__inv_2
X_6477_ _6475_/X _6796_/B vssd1 vssd1 vccd1 vccd1 _6766_/A sky130_fd_sc_hd__and2b_1
X_5428_ _5428_/A _5617_/A vssd1 vssd1 vccd1 vccd1 _6067_/A sky130_fd_sc_hd__and2_1
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5359_ _5359_/A _5461_/A vssd1 vssd1 vccd1 vccd1 _5360_/B sky130_fd_sc_hd__xnor2_1
XFILLER_101_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7029_ hold112/X _7018_/X _7028_/X _7021_/X vssd1 vssd1 vccd1 vccd1 _7189_/D sky130_fd_sc_hd__o211a_1
XFILLER_101_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7242__35 vssd1 vssd1 vccd1 vccd1 _7242__35/HI _7341_/A sky130_fd_sc_hd__conb_1
XFILLER_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4730_ _4730_/A _4730_/B vssd1 vssd1 vccd1 vccd1 _4731_/B sky130_fd_sc_hd__nor2_1
XFILLER_14_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4661_ _4733_/B _4660_/Y vssd1 vssd1 vccd1 vccd1 _4734_/A sky130_fd_sc_hd__nor2b_1
XFILLER_80_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7380_ _7380_/A _3670_/Y vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__ebufn_8
X_6400_ _6400_/A _6400_/B vssd1 vssd1 vccd1 vccd1 _6401_/B sky130_fd_sc_hd__xnor2_1
X_3612_ _3616_/A vssd1 vssd1 vccd1 vccd1 _3612_/Y sky130_fd_sc_hd__inv_2
X_4592_ hold70/A _6627_/A vssd1 vssd1 vccd1 vccd1 _4593_/B sky130_fd_sc_hd__and2_1
X_6331_ _6332_/A _6332_/B _6332_/C vssd1 vssd1 vccd1 vccd1 _6365_/A sky130_fd_sc_hd__o21a_1
XFILLER_88_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6262_ _6212_/A _6262_/B vssd1 vssd1 vccd1 vccd1 _6324_/A sky130_fd_sc_hd__and2b_1
X_5213_ _5213_/A _5213_/B vssd1 vssd1 vccd1 vccd1 _5215_/C sky130_fd_sc_hd__xnor2_1
X_6193_ _6102_/A _6102_/B _6192_/Y vssd1 vssd1 vccd1 vccd1 _6194_/B sky130_fd_sc_hd__a21oi_4
X_5144_ _5143_/X _4987_/A _4989_/B vssd1 vssd1 vccd1 vccd1 _5150_/A sky130_fd_sc_hd__a21o_1
X_5075_ _5075_/A _5117_/A vssd1 vssd1 vccd1 vccd1 _5093_/A sky130_fd_sc_hd__xnor2_1
X_4026_ _4026_/A _4026_/B vssd1 vssd1 vccd1 vccd1 _4039_/A sky130_fd_sc_hd__xor2_2
XFILLER_71_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5977_ _6659_/A _5986_/A vssd1 vssd1 vccd1 vccd1 _5978_/B sky130_fd_sc_hd__nand2_1
XFILLER_40_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4928_ _4928_/A _4928_/B vssd1 vssd1 vccd1 vccd1 _4932_/B sky130_fd_sc_hd__xnor2_1
XFILLER_100_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4859_ _6931_/A _5937_/B vssd1 vssd1 vccd1 vccd1 _4861_/B sky130_fd_sc_hd__xnor2_1
XFILLER_60_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6529_ _6529_/A _6529_/B vssd1 vssd1 vccd1 vccd1 _6539_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5900_ _5900_/A _5900_/B vssd1 vssd1 vccd1 vccd1 _5902_/B sky130_fd_sc_hd__or2_1
XFILLER_74_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6880_ _6879_/A _6877_/X _6878_/Y hold64/X vssd1 vssd1 vccd1 vccd1 hold66/A sky130_fd_sc_hd__o31a_1
X_5831_ _5833_/A _5833_/B vssd1 vssd1 vccd1 vccd1 _5871_/B sky130_fd_sc_hd__xnor2_1
XFILLER_61_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5762_ _5762_/A _5762_/B vssd1 vssd1 vccd1 vccd1 _5770_/A sky130_fd_sc_hd__xnor2_1
X_4713_ _4714_/A _4714_/B vssd1 vssd1 vccd1 vccd1 _4720_/B sky130_fd_sc_hd__xor2_1
X_5693_ _7023_/A _5873_/A vssd1 vssd1 vccd1 vccd1 _5723_/A sky130_fd_sc_hd__nand2_2
X_4644_ _4659_/A _4552_/C hold80/A vssd1 vssd1 vccd1 vccd1 _4645_/B sky130_fd_sc_hd__o21a_1
X_7432_ _7432_/A _3731_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[36] sky130_fd_sc_hd__ebufn_8
X_7363_ _7363_/A _3649_/Y vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__ebufn_8
X_4575_ _5597_/B _4844_/A _4744_/B vssd1 vssd1 vccd1 vccd1 _4668_/B sky130_fd_sc_hd__a21o_1
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6314_ _6314_/A _6314_/B vssd1 vssd1 vccd1 vccd1 _6314_/Y sky130_fd_sc_hd__nand2_1
XFILLER_89_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6245_ _6245_/A _6311_/B vssd1 vssd1 vccd1 vccd1 _6246_/B sky130_fd_sc_hd__xnor2_1
XFILLER_69_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6176_ _6301_/A _6794_/A _6850_/A vssd1 vssd1 vccd1 vccd1 _6245_/A sky130_fd_sc_hd__or3_2
XFILLER_84_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5127_ _5127_/A _5127_/B _5127_/C vssd1 vssd1 vccd1 vccd1 _5128_/B sky130_fd_sc_hd__nor3_1
XFILLER_84_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5058_ _7204_/Q vssd1 vssd1 vccd1 vccd1 hold87/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4009_ _4009_/A _4009_/B _5671_/B vssd1 vssd1 vccd1 vccd1 _4012_/A sky130_fd_sc_hd__and3_1
XFILLER_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_75_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold83 hold83/A vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_75_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_35_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_3 _5022_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4360_ _7070_/A _7202_/Q _5057_/B vssd1 vssd1 vccd1 vccd1 _4361_/B sky130_fd_sc_hd__o21a_1
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4291_ _4291_/A _4291_/B vssd1 vssd1 vccd1 vccd1 _4291_/X sky130_fd_sc_hd__and2_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7278__71 vssd1 vssd1 vccd1 vccd1 _7278__71/HI _7377_/A sky130_fd_sc_hd__conb_1
X_6030_ _6118_/A _6117_/B vssd1 vssd1 vccd1 vccd1 _6031_/B sky130_fd_sc_hd__nor2_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6932_ input3/X _7116_/B _6931_/Y _6846_/X vssd1 vssd1 vccd1 vccd1 _7154_/D sky130_fd_sc_hd__o211a_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6863_ _6875_/B _6863_/B vssd1 vssd1 vccd1 vccd1 _6873_/A sky130_fd_sc_hd__nand2_1
XFILLER_62_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5814_ _4465_/B _5812_/B _5839_/A vssd1 vssd1 vccd1 vccd1 _5849_/B sky130_fd_sc_hd__a21o_1
XFILLER_50_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6794_ _6794_/A _6794_/B vssd1 vssd1 vccd1 vccd1 _6865_/A sky130_fd_sc_hd__nand2_2
X_5745_ _5745_/A _5745_/B _5745_/C vssd1 vssd1 vccd1 vccd1 _5747_/A sky130_fd_sc_hd__or3_1
X_5676_ _5676_/A _6118_/A vssd1 vssd1 vccd1 vccd1 _6029_/B sky130_fd_sc_hd__or2_1
X_7415_ _7415_/A _3718_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[19] sky130_fd_sc_hd__ebufn_8
X_4627_ _4688_/A _4688_/B _4626_/X vssd1 vssd1 vccd1 vccd1 _4629_/B sky130_fd_sc_hd__a21oi_1
X_4558_ _4554_/A _4554_/B _4653_/A vssd1 vssd1 vccd1 vccd1 _4602_/B sky130_fd_sc_hd__o21ba_1
X_7346_ _7346_/A _3631_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[20] sky130_fd_sc_hd__ebufn_8
X_4489_ _4562_/A _4562_/B _4488_/Y vssd1 vssd1 vccd1 vccd1 _4523_/B sky130_fd_sc_hd__a21oi_2
XFILLER_77_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6228_ _6962_/A _6420_/B _6228_/C vssd1 vssd1 vccd1 vccd1 _6230_/A sky130_fd_sc_hd__and3_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6159_ _6524_/A _6966_/A vssd1 vssd1 vccd1 vccd1 _6160_/B sky130_fd_sc_hd__nor2_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3860_ _7198_/Q _7197_/Q vssd1 vssd1 vccd1 vccd1 _3861_/B sky130_fd_sc_hd__xor2_1
X_3791_ hold53/A _7202_/Q vssd1 vssd1 vccd1 vccd1 _4359_/B sky130_fd_sc_hd__xor2_2
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5530_ _5530_/A _5530_/B vssd1 vssd1 vccd1 vccd1 _5531_/C sky130_fd_sc_hd__xor2_1
XFILLER_31_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5461_ _5461_/A _5359_/A vssd1 vssd1 vccd1 vccd1 _5461_/X sky130_fd_sc_hd__or2b_1
X_4412_ _4412_/A _4412_/B vssd1 vssd1 vccd1 vccd1 _4541_/B sky130_fd_sc_hd__nor2_1
X_7200_ _7221_/CLK _7200_/D vssd1 vssd1 vccd1 vccd1 hold98/A sky130_fd_sc_hd__dfxtp_1
X_5392_ _5541_/B _5392_/B vssd1 vssd1 vccd1 vccd1 _5394_/C sky130_fd_sc_hd__or2_1
XFILLER_98_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4343_ _4236_/A _4236_/B _4342_/Y vssd1 vssd1 vccd1 vccd1 _4389_/A sky130_fd_sc_hd__o21ai_4
X_7131_ _7151_/CLK _7131_/D vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__dfxtp_1
XFILLER_98_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4274_ _7177_/Q vssd1 vssd1 vccd1 vccd1 _5734_/A sky130_fd_sc_hd__clkbuf_2
X_7062_ _7101_/A vssd1 vssd1 vccd1 vccd1 _7062_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6013_ _5594_/X hold28/X _5595_/X _6012_/X vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__o211a_1
XFILLER_39_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6915_ hold6/X _6893_/A _6914_/X vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__a21oi_1
XFILLER_82_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6846_ _7117_/A vssd1 vssd1 vccd1 vccd1 _6846_/X sky130_fd_sc_hd__clkbuf_4
X_6777_ _6777_/A _6777_/B vssd1 vssd1 vccd1 vccd1 _6792_/A sky130_fd_sc_hd__xnor2_1
XFILLER_50_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3989_ _7209_/Q _7196_/Q vssd1 vssd1 vccd1 vccd1 _4172_/B sky130_fd_sc_hd__xor2_2
X_5728_ _5727_/A _5728_/B vssd1 vssd1 vccd1 vccd1 _5728_/X sky130_fd_sc_hd__and2b_1
XFILLER_10_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5659_ _6466_/A _6439_/B _5692_/A vssd1 vssd1 vccd1 vccd1 _5682_/B sky130_fd_sc_hd__and3_1
X_7329_ _7329_/A _3740_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[3] sky130_fd_sc_hd__ebufn_8
XFILLER_2_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7248__41 vssd1 vssd1 vccd1 vccd1 _7248__41/HI _7347_/A sky130_fd_sc_hd__conb_1
XFILLER_49_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4961_ _5286_/A _5286_/B vssd1 vssd1 vccd1 vccd1 _5120_/B sky130_fd_sc_hd__xnor2_1
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4892_ _4892_/A _4892_/B vssd1 vssd1 vccd1 vccd1 _4899_/A sky130_fd_sc_hd__nand2_2
X_3912_ _3912_/A _3912_/B vssd1 vssd1 vccd1 vccd1 _3996_/A sky130_fd_sc_hd__xnor2_1
X_6700_ _6696_/X _6697_/Y _6699_/X vssd1 vssd1 vccd1 vccd1 _6700_/X sky130_fd_sc_hd__o21a_1
X_3843_ _7188_/Q _4506_/A vssd1 vssd1 vccd1 vccd1 _4009_/A sky130_fd_sc_hd__or2_1
X_6631_ _6631_/A _6631_/B vssd1 vssd1 vccd1 vccd1 _6653_/B sky130_fd_sc_hd__xnor2_1
XFILLER_32_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6562_ _6560_/A _6417_/B _6584_/B vssd1 vssd1 vccd1 vccd1 _6605_/A sky130_fd_sc_hd__a21oi_2
X_3774_ _7173_/Q vssd1 vssd1 vccd1 vccd1 _5615_/A sky130_fd_sc_hd__inv_2
X_6493_ _6938_/A _6507_/A _6493_/C vssd1 vssd1 vccd1 vccd1 _6493_/X sky130_fd_sc_hd__or3_1
X_5513_ _5513_/A _5513_/B _5513_/C vssd1 vssd1 vccd1 vccd1 _5514_/B sky130_fd_sc_hd__or3_1
X_5444_ _5444_/A _5444_/B vssd1 vssd1 vccd1 vccd1 _5445_/B sky130_fd_sc_hd__or2_1
XFILLER_99_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7114_ _7114_/A _7114_/B vssd1 vssd1 vccd1 vccd1 _7114_/X sky130_fd_sc_hd__or2_1
X_5375_ _5375_/A _5375_/B _5375_/C vssd1 vssd1 vccd1 vccd1 _5375_/X sky130_fd_sc_hd__and3_1
XFILLER_101_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4326_ _6761_/B _4326_/B vssd1 vssd1 vccd1 vccd1 _6421_/A sky130_fd_sc_hd__xnor2_4
XFILLER_101_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4257_ _4257_/A _4257_/B vssd1 vssd1 vccd1 vccd1 _4257_/X sky130_fd_sc_hd__or2_1
X_7045_ _7045_/A vssd1 vssd1 vccd1 vccd1 _7045_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_47_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4188_ _4188_/A _4188_/B vssd1 vssd1 vccd1 vccd1 _4238_/A sky130_fd_sc_hd__xnor2_1
XFILLER_55_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6829_ _6829_/A _6829_/B vssd1 vssd1 vccd1 vccd1 _6829_/Y sky130_fd_sc_hd__nand2_1
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5160_ _6240_/A _5611_/C vssd1 vssd1 vccd1 vccd1 _5161_/A sky130_fd_sc_hd__nand2_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5091_ _5091_/A _5091_/B vssd1 vssd1 vccd1 vccd1 _5092_/B sky130_fd_sc_hd__and2_1
X_4111_ _7181_/Q _7180_/Q vssd1 vssd1 vccd1 vccd1 _4377_/B sky130_fd_sc_hd__xor2_4
X_4042_ _4042_/A _4042_/B vssd1 vssd1 vccd1 vccd1 _4237_/B sky130_fd_sc_hd__xnor2_2
XFILLER_37_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5993_ _5987_/A _6577_/A _6674_/A vssd1 vssd1 vccd1 vccd1 _5993_/X sky130_fd_sc_hd__o21a_1
XFILLER_64_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4944_ hold75/A vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__inv_2
X_4875_ _7036_/A _7014_/A vssd1 vssd1 vccd1 vccd1 _4895_/B sky130_fd_sc_hd__nand2_2
XFILLER_32_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3826_ _7212_/Q _7199_/Q vssd1 vssd1 vccd1 vccd1 _3851_/B sky130_fd_sc_hd__xor2_1
X_6614_ _6241_/A _6613_/B _6704_/B vssd1 vssd1 vccd1 vccd1 _6619_/B sky130_fd_sc_hd__a21oi_1
X_3757_ _7169_/Q _7168_/Q vssd1 vssd1 vccd1 vccd1 _5625_/B sky130_fd_sc_hd__xor2_2
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6545_ _6546_/A _6546_/B vssd1 vssd1 vccd1 vccd1 _6547_/A sky130_fd_sc_hd__and2_1
X_3688_ _3691_/A vssd1 vssd1 vccd1 vccd1 _3688_/Y sky130_fd_sc_hd__inv_2
X_6476_ _6475_/B _6475_/C _6475_/D _6475_/A vssd1 vssd1 vccd1 vccd1 _6796_/B sky130_fd_sc_hd__a31o_1
X_5427_ _5615_/A _5895_/A vssd1 vssd1 vccd1 vccd1 _5617_/A sky130_fd_sc_hd__or2_1
XFILLER_58_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5358_ _5358_/A _5358_/B vssd1 vssd1 vccd1 vccd1 _5461_/A sky130_fd_sc_hd__xnor2_1
XFILLER_87_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4309_ _7178_/Q _7177_/Q vssd1 vssd1 vccd1 vccd1 _4745_/B sky130_fd_sc_hd__or2_1
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7028_ _7028_/A _7038_/B vssd1 vssd1 vccd1 vccd1 _7028_/X sky130_fd_sc_hd__or2_1
XFILLER_28_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5289_ _5289_/A _5289_/B _5289_/C vssd1 vssd1 vccd1 vccd1 _5290_/B sky130_fd_sc_hd__and3_1
XFILLER_101_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4660_ _6475_/A _4660_/B vssd1 vssd1 vccd1 vccd1 _4660_/Y sky130_fd_sc_hd__xnor2_1
X_3611_ _3742_/A vssd1 vssd1 vccd1 vccd1 _3616_/A sky130_fd_sc_hd__buf_8
X_4591_ _5619_/B vssd1 vssd1 vccd1 vccd1 _6627_/A sky130_fd_sc_hd__buf_2
X_6330_ _6330_/A _6330_/B vssd1 vssd1 vccd1 vccd1 _6332_/C sky130_fd_sc_hd__and2_1
X_6261_ _6261_/A vssd1 vssd1 vccd1 vccd1 _6261_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5212_ _5210_/Y _5335_/B hold84/A _5210_/A vssd1 vssd1 vccd1 vccd1 _5213_/B sky130_fd_sc_hd__o2bb2a_1
X_6192_ _6192_/A _6192_/B vssd1 vssd1 vccd1 vccd1 _6192_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5143_ _6455_/A vssd1 vssd1 vccd1 vccd1 _5143_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_96_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5074_ _4366_/A _4366_/B _5073_/Y vssd1 vssd1 vccd1 vccd1 _5117_/A sky130_fd_sc_hd__a21oi_1
X_4025_ _4025_/A _4025_/B vssd1 vssd1 vccd1 vccd1 _4120_/A sky130_fd_sc_hd__xnor2_2
XFILLER_71_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5976_ _6997_/A _5985_/B vssd1 vssd1 vccd1 vccd1 _5986_/A sky130_fd_sc_hd__nand2_1
XFILLER_52_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4927_ _4927_/A _4927_/B vssd1 vssd1 vccd1 vccd1 _4928_/B sky130_fd_sc_hd__nor2_1
XFILLER_33_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4858_ _4858_/A _4858_/B _4895_/A vssd1 vssd1 vccd1 vccd1 _4878_/A sky130_fd_sc_hd__or3_2
XFILLER_20_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3809_ _4477_/A _4477_/B vssd1 vssd1 vccd1 vccd1 _4633_/A sky130_fd_sc_hd__nor2_1
X_4789_ hold97/A _4789_/B vssd1 vssd1 vccd1 vccd1 _4864_/A sky130_fd_sc_hd__xor2_1
X_6528_ _6528_/A _6528_/B vssd1 vssd1 vccd1 vccd1 _6552_/B sky130_fd_sc_hd__or2_1
X_6459_ _6728_/A _6459_/B vssd1 vssd1 vccd1 vccd1 _6461_/A sky130_fd_sc_hd__nor2_1
XFILLER_69_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7302__95 vssd1 vssd1 vccd1 vccd1 _7302__95/HI _7410_/A sky130_fd_sc_hd__conb_1
XFILLER_48_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5830_ _5872_/A _5872_/B _5829_/X vssd1 vssd1 vccd1 vccd1 _5833_/B sky130_fd_sc_hd__a21oi_1
XFILLER_22_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5761_ _5774_/A vssd1 vssd1 vccd1 vccd1 _5761_/Y sky130_fd_sc_hd__inv_2
X_4712_ _4756_/A _4756_/B _4711_/X vssd1 vssd1 vccd1 vccd1 _4714_/B sky130_fd_sc_hd__a21oi_1
X_5692_ _5692_/A _5721_/A vssd1 vssd1 vccd1 vccd1 _5696_/A sky130_fd_sc_hd__xnor2_4
X_7431_ _7431_/A _3730_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[35] sky130_fd_sc_hd__ebufn_8
X_4643_ _4650_/A _4650_/B vssd1 vssd1 vccd1 vccd1 _4655_/A sky130_fd_sc_hd__nand2_1
X_4574_ _4744_/B _5850_/B vssd1 vssd1 vccd1 vccd1 _4844_/A sky130_fd_sc_hd__nor2_1
X_7362_ _7362_/A _3647_/Y vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_hd__ebufn_8
X_6313_ _6313_/A _6313_/B vssd1 vssd1 vccd1 vccd1 _6316_/A sky130_fd_sc_hd__xnor2_2
X_6244_ _6244_/A _6244_/B vssd1 vssd1 vccd1 vccd1 _6311_/B sky130_fd_sc_hd__xnor2_1
XFILLER_39_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6175_ _6956_/A _6160_/B _6962_/A vssd1 vssd1 vccd1 vccd1 _6177_/A sky130_fd_sc_hd__o21a_1
XFILLER_84_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5126_ _5127_/A _5127_/B _5127_/C vssd1 vssd1 vccd1 vccd1 _5284_/A sky130_fd_sc_hd__o21a_1
XFILLER_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5057_ _5062_/C _5057_/B vssd1 vssd1 vccd1 vccd1 _5203_/A sky130_fd_sc_hd__nor2_1
X_4008_ _4008_/A _4008_/B vssd1 vssd1 vccd1 vccd1 _4016_/A sky130_fd_sc_hd__xnor2_1
XFILLER_53_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5959_ _6674_/A vssd1 vssd1 vccd1 vccd1 _6665_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_48_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__clkbuf_2
XFILLER_45_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_4 _6956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4290_ _4291_/A _4291_/B vssd1 vssd1 vccd1 vccd1 _4334_/B sky130_fd_sc_hd__xor2_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7293__86 vssd1 vssd1 vccd1 vccd1 _7293__86/HI _7401_/A sky130_fd_sc_hd__conb_1
XFILLER_27_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6931_ _6931_/A _6933_/B vssd1 vssd1 vccd1 vccd1 _6931_/Y sky130_fd_sc_hd__nand2_1
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6862_ _6862_/A _6862_/B _6862_/C vssd1 vssd1 vccd1 vccd1 _6863_/B sky130_fd_sc_hd__or3_1
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5813_ _5838_/B _5813_/B vssd1 vssd1 vccd1 vccd1 _5839_/A sky130_fd_sc_hd__and2b_1
X_6793_ _6793_/A _6793_/B vssd1 vssd1 vccd1 vccd1 _6814_/B sky130_fd_sc_hd__nand2_1
X_5744_ _5744_/A _5744_/B vssd1 vssd1 vccd1 vccd1 _5745_/C sky130_fd_sc_hd__xor2_1
X_5675_ _5674_/B _7190_/Q vssd1 vssd1 vccd1 vccd1 _6118_/A sky130_fd_sc_hd__and2b_1
X_7414_ _7414_/A _3720_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[18] sky130_fd_sc_hd__ebufn_8
X_4626_ _4625_/A _4626_/B vssd1 vssd1 vccd1 vccd1 _4626_/X sky130_fd_sc_hd__and2b_1
X_7345_ _7345_/A _3629_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[19] sky130_fd_sc_hd__ebufn_8
X_4557_ _4652_/A _4652_/B vssd1 vssd1 vccd1 vccd1 _4653_/A sky130_fd_sc_hd__nor2_1
X_4488_ _4488_/A _4488_/B vssd1 vssd1 vccd1 vccd1 _4488_/Y sky130_fd_sc_hd__nor2_1
XFILLER_1_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6227_ _6537_/B vssd1 vssd1 vccd1 vccd1 _6420_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6158_ _6528_/A _6301_/A vssd1 vssd1 vccd1 vccd1 _6158_/Y sky130_fd_sc_hd__nor2_1
XFILLER_85_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5109_ _4632_/A _4632_/B _5108_/X vssd1 vssd1 vccd1 vccd1 _5116_/B sky130_fd_sc_hd__a21o_2
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6089_ _6089_/A _6089_/B vssd1 vssd1 vccd1 vccd1 _6186_/A sky130_fd_sc_hd__xnor2_2
XFILLER_57_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3790_ hold58/A _5056_/B vssd1 vssd1 vccd1 vccd1 _4355_/A sky130_fd_sc_hd__or2_1
XFILLER_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5460_ _5521_/A _5521_/B vssd1 vssd1 vccd1 vccd1 _5463_/A sky130_fd_sc_hd__xnor2_1
X_4411_ _4411_/A vssd1 vssd1 vccd1 vccd1 _7085_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_99_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5391_ _5391_/A _5391_/B _6455_/A vssd1 vssd1 vccd1 vccd1 _5392_/B sky130_fd_sc_hd__and3_1
X_4342_ _4342_/A _4342_/B vssd1 vssd1 vccd1 vccd1 _4342_/Y sky130_fd_sc_hd__nand2_1
X_7130_ _7151_/CLK _7130_/D vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__dfxtp_1
XFILLER_98_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7061_ hold127/X _7045_/X _7059_/X _7060_/X vssd1 vssd1 vccd1 vccd1 _7201_/D sky130_fd_sc_hd__o211a_1
X_4273_ _4379_/A _4315_/B _4272_/X vssd1 vssd1 vccd1 vccd1 _4334_/A sky130_fd_sc_hd__o21ai_1
XFILLER_86_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6012_ _6010_/X _6011_/Y hold63/A vssd1 vssd1 vccd1 vccd1 _6012_/X sky130_fd_sc_hd__a21o_2
.ends

